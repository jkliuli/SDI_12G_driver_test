`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
HaBQz1qtMJbx283nr4KZ/krD+gxavgbulj/CM6g/uFii/Hf3PR0pozrRlLLErcbE
T9PIRF53Q9WBauSKtlcu1qBS9CEM9vPyUqKTKzc/WIoFj5pByIYDjZGNd1BCqoQ7
sUP4cznVzEY/XrS0Jd9f5PeYI5W6dG/rVOpnRrPX8VQ=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4080), data_block
tm15BEpytGQ7XCqeeYuoilWqL0gNd7pEmNoPQ+gBCEZPs7ZZWICTeRxaXNzgWOsI
Y5GO36+Y05HrUl0jDBkMMpFamqsUIjl6u0b7Hn6CviGe+tpnPDaLPTbSAsldUnjw
nijgW5dJiOXgwqBp+t4DxyUOrpBLMU82Rp/DlENQ8rTFMEm1bk2tDY1yiRJA1H2C
Bi12Ief+xRjo/aCzUvyI+qsLF1ICg0ZDmVsvtvSxx66YULMPyeYjulIYhC+URlTa
5PZRe5OZGc79lwU8HrJkR46YgUaxcxCAMjOMEfL4gu4yZG43thEQQJxW6k1pBmB4
JmElvrTQ5a9S6GCYFbRL2OLSYm1eWsybKiP4WcJcRQ3zVocUNkKfIgNxRPLmtCco
/TSviGYA6fLCO3SbYa199Ju6o7aRfk0DbtJ4cOx77iFgJYYX87eUDCI46xftFxiz
Itt/IaAA4vp4I+yLvdzUPlSihzEw460zwoiUsXPlXQ6rMI6qSJ64A+aWBEeWX5vZ
GCWe3DXuPjK4/ukUmcfG7Pj2SEZGwyiY1o+S3zvB/SAe+dBdMYWRETQaGrXk0cCw
f/PBYKI6dPQcN8nAEq/m1MHhHVg8ZHqKY6BAJ4HIRzxVqFT6RZeNSD9yr29Gbn/f
1tFvf1KMQ82i/cTuYjZWA0VC8oQBiuFDtQwNNRKqoHONRi4DSRVKtu8QZFywcBgP
ml+xGyMlyra4/L5AnR64r5Y4xejzua3Jm49YNSljc534T9QmyjTIJY8NMSFuN/+w
/sM0/pXdw4jqQN4wvYva75sRojLPA0TF2Vyi/fmUmsqesxXc5NjmIAgHYgi47HtS
sw9qoZejJsC15YURlPDSD91EXRTmqUm9OhNVQf4kkK3YMwJJp8nSa82np+MeDMNO
M191Y6i3/niF6WYF6nvTtT7AlJfPjjrKDrugy9MfCLf2ReVWBZUpentpEB3Drpnt
5ANu7mB0OS3OxdhZSQ3AjtyIVn0Wt5Wy6LXbyEM4nIdO6c5CBWD5ACpVxb+U7upV
ixM1qFYuMWHnzXRYxnJ3cfQg8fUMp8RcaT51hhvFYheKvqFZj6Mm9bkGW8KlDTE3
2C8coWSNl4wndhjtT9xBIwL52aYr8QYDfdfSDV4ZYqRTmpMOh7IKPMZM67KyLIvj
+4zxWRupF9dUT6smDsxh1yPbmLzqlrfFHdUam5hHecN1y25u+muxwvkkIlzclRq1
Gf3HI1EOGORD/N9LWWws3DfgnTk2dl8ZKS2zOME8eejzelgr0CFk+4qPIRCoKYAM
vyJzzV8tORVhkagn3T2qg8T02hC0MPaoGMjTAglzr3a0OPk4e1PZQiaIq2HT8bEp
zFZw3wFSViQb8Uyky6VbpoYCjiQ4OMN8t8hyA4uv2NVmsSP/wfvNT7BGtmOLBJaA
lqolZwv8mJeh3FVvYJBID6hhTfc/aRhvtzlMmM/CYpTKargqxTeyT+67x4fqEAWZ
fLRIc6U+TZIiDWOGO4FXa+qjQtPoYKOkX+63z+48K965zYbJXawPN+FEhJkJyKAQ
lv3J7AvYEKm9cJcWhn3OcC70LkCqM2t/6LgSbqiMpdJyKPX5EhtMC5MqbJFXwiv6
ynJrI6Ue+fa6P5uT4yeVc/GUbxSzWMxiP1iazvuqvnCAXknV3aezw+S4olAIHYRg
oRKbQKjUv3snlrYMVwPPkJdEbaOzdxwKAVPWnPwKxbnuIdgWe95oEcW9gj7HiKik
5CjANsischW8rBRVO+7QeRnblZoiMB8mV4dcMdr8zFC6Ezi7iM+CAtIR5w2GdkGQ
X0UmphMwIlx/If8+q/A6D6q45OxsfWxJ2TfJVHq6sKnp60d4anP8XByMluYZxbT9
gNXJdCb8M5yTjracMVy+i0q0pWrCCGnAsSRT8EneFRfm0Gx+EksPcGhsMQWJUC5P
rnwM3rLNGguZ435nQ5xav0e9KGeGdwbropZhTD3w9dRucYYZjKJt+8Tr/MuuNl3J
h4885ITeaD8Y1VcY7o/YJSUQJoiWixvgdAZV52fe8GiLi3BSOyQDXAa2HmaQMnzj
uKbbRjCKSVpR+pnSqJJsi+dZkwIwShFjgCE4Au/FiROSfTARFGFThLmnMeItmAMh
v1qS/lS6W3iKGkYDCqg96zsc+ETdepOSEXNLBc1xTJXmwK5NixDiB67cy4I2d8EM
uxRX5lk+lVRLXBvBa+7+7DmncKQ2vswxp27kXljkU4RQFS2Mr5mrezxqn+dXi+n0
eBZT3kuyDd8vQ8i7E8gJsKF+f52n7sdsp9LPGndd4NlPlR4sy+4TulbFxXgtEle1
baZSgWD02Mb8je2DqJko2o4HkX91Mv+Rf3PfW/LkXqrKppd4sCMd/ALgJnopAMLq
6tnkPLgiuN0GEJllD4sovQMznjocbPWuP3uVwbiZ20hsnOldMfUGSbOurYTz5NOV
TIQS57IG6eN2eN6EC+vVuxKji5ly5ow9ot8ONG5CLTw9dPASzqgCKavswWESYdp0
p4cVsRLh8ryvjMehwix2gA01EfJPfxuA2xhVsnxe3dIvCKIi164ImRzw58nY6QwC
Ojt86v+Q+8A7PEYvbgeGF9bY7HGDJwNTTzc82wVQ0RRiwaP13RNmU6Jil1loTOUX
XV3EBWU2APDSwRVW8Ce22eeb1i3dqYTrqyOM188iUlg1HbELOwrHDPKgSUsd1UaP
LH+xwD+woLr10cNGutKj+MGMug78Fpr4MPo6jUe+9us8IswFbnvMNXmTNvF9KRLS
a07aVqx4q2x1/6oIAWciaLLfG894OjeV3igCZyAueMKLkRYNEK3q3wsQipsxHV6K
yliqAMkdnvHE+D53mDoTRYaXedHPkddu4IKKIef5eGCQjT7hR5wl6Ujyx4xhd3zw
CmWORjbfWjyMR5o8KSUTa1L7UOF3HciaBO/vY6Os6F8TDoryrQ0wUilA+TShRQ+B
a6kVHCcpQsqd35KJN1PvKAJl250RqsqMH+FidjwhWjNvwOUvG6JkJ1we+lMfB3EI
IL3w5cGWP6F0Eqysaib3PmU4NWBaGSYnCoFnC9oguEKC0c0JL+vAlHhdjjW4gA+6
9hlm8qYHCJ3qMxgUuPn3XPPhwA+nNSbMdKU3Vpkt5PdGvCkY9fApb6itqHlWreZ2
IvoYNVELHggFVsiS1xszWI8IWlZi+vPnkxXKcbqKF7Tur2EyWL22GopKlPPaV2rs
UYc47Cp8bxPf8jPcGZ3wVLH47DS0ucaZ7s8+dvdll8kVv56odKvOctJDmqGh1THO
v17sOhidI7Xp073I38f7qxISgZSxWeagXolxWfd2dPVLXXDrguJ317pyNgAa+MM+
KWfLxGasrkZiLkfHQDxUhcs9wnyAj+60HQWXl2jgDMFtJaFhU+t/DKk1q3OgCspe
f83G+Z3G/CO4YNbgvpnb2T6+Vq4rHwzog6F0UJUwtxeaEQ1XHHWsPrFutwV2nmY6
1DlI0Hqjdpp8I4jQ+6tjL9gw/278Zq0BEb/lZLpV9+JhXsXbBi1yENt7lysHQIvo
4/1sdt1PoUmweFjmr84tzGqPLJaqImZUJHVTWp+2GeJ7WO4V4LYcUx3sVfrCd5s0
g1H6TwXXmN3M+kLQeD7aDJE7CpRTUSWxOxc7X88G/45Mbtmq8Ogk36FWd/CVlGxa
soOz4BemjjTQMEK8zMJsxbJXs/cnLpJqjVeaVgMWnQLwEdu/ZOhFoA8bl+GTJ5EX
gMgAlX37tucPgCQ1cBe5GL6D0gD83mzovdLnVGVxbge8r6Vj+H1YqbY1jbb8aNgj
X/rj6lFc5Jq94XWYTGBpJg9oPRMoT6guylbfVz3FlpE+U4En9Q7453j6QGMyJlQu
v9iGA7i5+HODf5fDMDm+Dn1kmfN2r88fzAFXWSdvtSbMoiYyMEbURxh6oIutZhOO
6/nKnRX+z4D7qkLqGAZT+5+gJzPLO4G3l8jMvK2KnyboKHEHkMZxFylctwQ1P8Fh
CD8Bi79YSgINN/m9aVnWT4i5JOe8Wy68sH20D6zguW33nWOuL81N2judaboWhPFJ
ebQHVnjPeBi1rF2I1YaOlwpMkjKLZjy8fOS0ygnLIAj+pBMTLgdI8GlxDYVBVfSR
7rhPFWf+gAAEJahRREjsHcV0Of0l3Bb4BP+i5GlNMDlcyrjCeBlov4fbkQRwyylT
mJ4U0rWeIVlFeFbWDv1+YwBsH+0cUcHi7a0p0uLCbZgYkGI5JQY+SMh+IgwoHHV0
5/kVlhJhhW04Cg+NwrZ6Fkz8LgZrrjkg6GGdshMRXZ3K3mCTKGZvRnEpF1tOfjE7
i5ddcnGOCqBKyCFpaeC3zc4qrI6GtfwOZbQ42i3kLHyfLkDq2mrfzFmjDK+sk+I/
o5dvvUzuR1Jk5LGxMhkrA7C8eLLjjDAEvsPJqo84ldRKxW6l3Qc2GPzFfj9t3UAj
GmbAYuiOGQIbBdeZDvx7MzSZRYHrPCmLMwRpyyhICXQBG9LUAvs7W/zpjd1PNaQo
IMaUWSzWARU13s0ORCEzBTyPdEI0quO3b5IyroyCHurituhOxgRPV3OsGypt71Nu
CY7ld/m/TROYbP1UkikjQJYZ08Mi4cBzb4qJc/NygnH5H/jzISAW0XND7FGHNPFf
H2XQV5fxTCe/JzboEYX7mzJenh3Iym+6sJuKi7axA/LkqisIrDYP1RElIy6E7+Lj
dwn71xvByPYZSkQMZPX9aen2IQXiMypMH/UETbuJrIT3kPfObxeXL2qlHA+J4Tbz
0ROGMW3T1mwDovxGeWwMsR3idjqYImmz91pf2YZE3p0wbzs0ejivC6WZyAOQcK7T
Dz3oqUIFZ5f7JR+5Y+yAsk8VxwANT41K2lH26FVSD5sBxXBfQwgr1kyOSQIuHZz3
3icNnVUif8j/gzGFFyd/REyi0fkkwK9E9ohD2AmHzkI3Wv4VdjI3NuJPR7EFq6rS
CQClV0PKs30QFUK0w2ZbthQszGxAZ3E94Jnc9plOgA2knhF0aqEL3jb/dQpfkE/E
4rZTuSgC3ZeOMlj9I2rdzD4IGjUe5tJOKBtpBTjtMjsLQOYzVCi5ui181RO1fyF2
eDKuxjSfGso7WGr8lK83k6LJ/JfrtZD7jpA+S00eLqDtqkiSaJbfXaxXAf/wLqwa
PvczW56NA0ho1G1+Xf4Ddmj0x1KYYS3OnAWffPOVELlXuKLuZQg8tHEN5tQgMOqX
WFbwhp39Y+j68HQcYWbH9hOdA8eYgHygJGGRMlPCiO3kmcSeoWlPmHLJUqZJMVW5
V35+NYzBQzWLvSKk6+qixBwi+DwsT6OTAZil3ZVG6z9EQTtzSZ6zC83T+mI6dmW+
zdaKzQHtqhmd2QiW6xdMXAm31GH3+tvDEAIMUu47yPbAGBH7snEw3uXEt7bdpQOw
JRO8feQreuBRK1N5ETDt8yELfrUBavRKYx+8nfSE1NtzwwL/VusKxnmacW9mUwnN
`pragma protect end_protected
