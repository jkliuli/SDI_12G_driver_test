`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
ez3nirT/g0facimvB+0D+3HRBoVBkIKwBGi+DtDS7BmY00FBT1HEP/bhisGyufAP
GppEJghRZjLByBr1BrbLuSz6Yuo+gDEqifEk05Xy7Qg5+jPEq0eE5SkQccexKEeR
Ik7mClukymC6iVm5QNSP9OnR5QmxhbMjk4i8DvTQxvs=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 31712), data_block
CbBDIVhRNTd98YeBesKcwdV61YyZkUZZSiHwxmD5APobOzLq/GAAk4hJv7lsytON
SpCH9Zl/UjBhURVlE8aM9ZRCB62SgriKn17I2zATessrplnuWwbpvRgQsokxMln5
MqPHHF32OkWxPxgVTkytzlUysKJpO8Thc8YhuMlzTHS8gSgywDNVVFnjXWPG+XjO
2m8r+vFvpssurOogK0k0zCkm5Sazm9nnKMWtnbgeplYvkVaQzc6NNNYexUZC3jRW
Fm+IqhPqRT22pWY4FiUbQtcF3FsKMVfmFxJHQx2wGBb7N08G3uU2LfP/yULn1z8n
AVvEmDJg7aGhW/O14SQk5SQXewl4yhG8Csqx8j3mhXl+rCPTrSz1kqa77xU7Bl63
umIMR0jHugCkA7aivvkxsaPgMdV33BPyMVkPQHX8duIHxeSWouHVJJx8EhKmBkzd
S4PbigdJ5JtHpwjUWK4+UoRUjP8Ur/7fvMMB60WoqhX7ysYH/BhqRvTrB5sQqEHw
si3aOpRv7mqWyKnU4Pn9gQt/k37u7ufBPpfhpDjyj/li4TH4l8NQXj9gWplp294x
YvB4Iw/aNOag4FIxnTXWz8ckIWQJJLNqE/z7SuDZDlbqrOp8NyMEc8dtSTuIFIt/
3EnlzaKU3tffsic+OY2iM/MmUJuoeFts2o9FcCookp82ep2f1KPTeVzTzXa4o07u
KfyvQh+PG6xJQQzLu0eibS0lEtBKT6A+bq7bMFtub9bndyp+to4Z7p4ODpCg9QkH
ZJD8G+/X0gJrEireDBCm8ZnGQw7hVX3V20sQkiyKfy/u6HaxhAsR1WYuMp6Yj4yE
3GXwEknD8G/bZDFBfXidnPNOyuGR+kOGee0dfy28XqEOERryBLapPVNE3PmHImo3
Bo+o2XN4VneryZKnK7YIYeHbEpao2WRvcg0hg29BZNER5SDVTGaFE2QAdYCDweSB
Ti9dL8lFo/TrD/v1ywk7MGq9MGYbYyuExS7I64+PYqk/DXQS2ZDO5khMheAkbTiw
HG3ZTTw9S6pppBLPCD0PpAteCzJhaiSpR/YrUoQ2uGPnKPju3Ik3XW9jGhGPwZPJ
RGzPQfsmKJhBlBRqoeNEdpNDCboqVgTp7coATy0JiGkcLZMoI3nc3BHSif7oib0J
Tp5MAcyeAsJdgMe7ky2hv+fWCQkQZisd4J8a1nt76b/s4xy+xReGNUVObubim4zg
FLu6mr828QqTrAncEyiJfQ34c4AvRVD5V3JEmT2MrD2NmibSaqydPmhFriVcL0gq
4rKV1dXfN4M25but+4PNFGHdknZxkEkHlTtmwMqzECmh51AKk1oW+X5UrbPIvY4K
391NhD/EmX8XpcXfmIe7G4uevlWKnuYEjBIyRlHpXwLeRlIbt+E8nL8LEU5cYTzD
78G1XUmV3F86R4RIfObPboD2uZ9Z7f8zDm5qfZmcExPd1vjYx+GD3AaXKYIB4XSA
EAxIicFFmemre2SZWFVCDX7nIhZRibFuZoDhYbaXQc74HfGLhSdJV5mR/SeBv++C
KqBQSRPlpuebNl2SfopOOTa26RLgrFlmGeTsAJimrF3perGCJeylUooNUmInyfz/
SPCV9d7dNbVJeeLvmrvUgTVPV+l/DzyldQ3gSeD/a0nfXTZGvYXhF9ZDLS0CbsS4
WQS4QU68TmIu27VSpoPuZTAI/rzFxswZhicXK7J7xTxvJ/rZDDvfIbaYAG6IJ/Lq
1Omiyq8Ay/eU26plJqrYVCHZQtaP2i2QKJp88bKOsYFKgnmZ3cTM6fYEZeDIMY9h
zcWxjy5g+SF0MbCwkwwGJVB3TMOwJhEmIuZ+O2+axSSVlj4fLz6pS9xJUUnl+qpR
EV2cUA5634DWd/jgEn0A3bLOyzO2Xwf3q5aoLNnaOrNgdj8AKYOG+GHJM663HZnj
uVPLn34fo/tFXWxFoc+ivK5cA9aNRtJUG7YsjWb9Tv3cBkVTx/pSmN6OHaCpEz4f
vEbyVv9sJceyMEGJsSfzVW3f2FHFN+FM9aeQxJCAmJxFkliCTKCQ0Y8ENWBdFAUc
sd4BfQh1n7cbUG1RJUcggo0WpTLIUZNAhTtms2gaqQJfmRIGt6o6Mx1Lo3rg1Esh
Gc7KTH9gXWQfCVOP9HVeKvJK+BAY/aurS8p1kRlBgUuNR2FWFzJ2d91u9ngMoaH0
K4Nn3MUaUh7Q/kbO7MQEbb8sOw/9R1thsoE4w0qqPzP2D8V8Cobef8/KmfQWs/vr
+q3RPM7+jwlvmmW/HEBSJQ6xCiuPQ1Punk6ZZzASgMkrBRtp663w8D35kTl8hxar
sdQgGa3DiDmH8B2/splgN5QOFA7A7IqE1go+Wic9/MKcy7mtFPCkI0keKrXHqJ+S
fp12jSACBYp79WPhiyy8J6SuP5rrlL2IZrMbcMmPlsHN+eTV7jlSLhnNLpvUwnRX
lSlrQLQpK1/56/X4go8TTFE5JwSBylQ41Cple0subRdxQT/B18hbWiCVZxPHgivl
sacaYYpt1MbHu7iKWGaDsHaFk4CBByc1pq+zQwBczDFCIFSi6sWVUFu4rWF9DG9c
IrMd44GII4PV5uKaDAznMt4ht1VNDU/5Ykvu2KhPGTLNV+uZif0Fma9t1zfWQiMl
rZU94OqAVYvfzIkSCAycWjj16TLEeoTLE4L5l+qCWSWVj9L0TyUqQncUdXgA2dVr
xIin5VRbQVbQPVx0USOUfOxwZDBUOpCe+rNSXIAg9GlSc2J0cifkkHF4X2gZ2mYf
YOd8WNCKCqenaJBi8jFlnBcLKyx/kXpnmVpgswwPNfk6+qkIdUaUptFPIjT0SGhD
gDTRYM60mK/YlyqIUA48C/yvXAS5SJmRGNKn/MlWpBqHWVxL95DSEq7FA2fkGQDo
/KK+2nau7jIZnPWag0ixroxV1u6lKP7JSq+QWh8Ro+nIIz2qJdxWtqfLyVcJnAl+
PAvGxU96QtJJcB4CPgxQfzq6Yz/Hti8rvyVF1rYa9vZI4U3wArU7q1vyq43l3dfa
s0meTa4ddKsnAT9uHIwjhwcOJP4QhZ6TaE5M4ylFVRlmKDMEI0nlWjdAIqDDjfmf
lz9ZBEhy+gjbEBLsIC178MthfNVWV2jC2vLg1UMcQyzxVunHWZWcUgGc1Dc/BmZR
wAONTPqlJycR6/bZNb8yNH2NEr/rt3K49qqOFpD+3/wVpj68Mpmcj7W7rlC9aaBn
a9FF4iEf69D34b+krRY1osLcG+59oFtle2gsgk+S4EXUomedgwNMZlORacoEGwFF
xQSuStEvzZMT2orsGGVZYiF9iZwjBIod8DcJlC18Wreu0bJZqQjI2xjp9fSv7GWu
8g0tZmWNlTMIeBjaqD/6ljnazCA4pTtLxwgyHRz/FZnHtt5VO2d1Rba6x02v7mB0
Wg+78phOC5iGYm4IX3Pfr2yTpp7oU1TKSZSvwNQB0oAL30/H5mcVfCmgUyjIEJ6c
8De6MZ5ub21fO12uPwAekV2sdIHmvQLeZ0zg+gE4tdGbjiMQPtLp2jRHQosiRb0/
C6Z9tYBiiT1v47sOzqjMGVa2Bqsb3/RgUo3gdMXuyyWQ9PUwD0LAsRrUrpJ1LUtB
IiphiT0XkCcEbxmJw5C6+4VVkBSk7tUVnzLQ6kRNqtPTB0ZiSeIqMYyoSrMzn6cW
ZMQBkf8/dKgwq0XvzICagE4eQ6G+Kgewtg33XHWM1ws8Exky6w0MnOlE9EZpZy1U
TfnggduUnyhrCBtkJyZ+hPJX/kqMyIrFwQLu/zM/NJHWAUQ5ibZstbx68eddW7zC
cHgufOteOOLYj8B8cTqB5fUTeDQsuZb+HDoHJJDUGmW7Lyp/myAXQ6tW2d4+Efb6
ISRvWNjrqgtej1UXh69Inw1KkDIgZ9sdJhZdQ1/oOxJMcLPEhC82atWMXtCQ7pPs
7Biw2ykFohDRPZRE252kIyfITjpcgegkZM58/q6RBrBTfkWQRAVHWTuK+O1RPeAt
JRPUax8+OpNhwMzteCHmy2nEpNaUYqVDT/gEywSlO6qW2UXMdHQ2tZy/YLWFhnA+
0e99qJTk7/AMwOguksuQ5IML+yk7F/1avryDSdiefhor1Z9nNAulxp8qDyRF0VN7
cSpc5djTMOfGFyrQnEiHU6vfKfoLr0EWMuYxITlohL6VEi7dCsZBGdSvY1zRFM5d
8Hx+gUy6/5CAVJ3SQqIjIEyYTw4AVpWL4EkRWshBVo9BLYHUjrulpZGyC7atAQUX
aq3BfapXMLRQn/lz3Zq8hWiTzLoqJualcgO8pCU8zBlMwK3bAbz9F+A5I2mwuzTK
iV+3sGz7c2TRBoYDiqVBEgU0Pgx2X0fcUeV0Aws5yhIWaC5lSCgngAR9xhnoj0aT
lCby1wY6Jg5vFcGT4BvWiS4UzmkAvr+WPKL93Qpg7jwnTXuhykzc579DKd8IcvMs
4aI93g2o2wiAP3ruImfGiiHazlkU7x9vVH+EfoV1q3+xDAGa5n43/rBqQpsni2E/
cm5ge2eUjh2yB5TFGPHEzawWBOwyOG0HQ3zWwoyzqaqYPWiUM0VdKUPTSjqDTU62
pmN/79VhWprFlv+ufJ44nfkqZb7nl6zK3GboYvV5kpxeMwMNDARVyb9QGwZAIRHw
mnq4x0xRPXpjEclsZ3k6FtZo0wxmHjQbVUjv/2gHRKBpLwofrUqtRLQEzHHT6csd
QQvpdjLwQY6FX+lVMs07lkiXB5Otqa1QS1bVM4I1LTSdoyXFQYu/QP8w5LWtfnB9
i7G6Ygd6Jcd4VQTT09xfziR+BPs6OfK0ohJ50QaoJ0i19DtQluLFjwOouy3xvmYW
FLmilvJV1TPK1x2QYjVH6CyXH0XOT/rJQrWWdzsZel5roYDwo5V8YXlcqahdZoTn
uROpRPnlx1e1cWk01SZe12e1Fj92oui2s2YgHobwvlDIQS6zux16B5Znx9wX6wzR
YGMf/p0LL/Xh/8xptWmXsSUj4Jt/8GQq0zvu0QOSdb5T7MEB+Uo9SxK3nRiRxjUg
FPTIGzeim5Y6s7Ajt32QIj4peHEnYsBKJhrz7U6pk5K0nmp43MUhmiFOq6IHdYlN
Jlh6hDzGQ0blazPigqR9lZzaizkUhomU30hXK0RpH2OfEWF+r+kDrTRcjpTaWnuZ
g/G/8hcFevaLX2Wn1GX1t31xVgzDP2nes7xJstsDhy5Ewd5KrWBjmyaZc4NGt8HI
LsaHOUj7aDXHyPioRl32eGRbbJl2QEkEHr1UExkwDPAljwiSGjQVQnOo9E+rDR53
ZYAc1OqF+HnVJdYvhmcnFCVmjj/i8JHpYCUFSAiXBxWxKNssc0L2W9g6gzwOHa81
1YrcrXRUBifJh54cvEby4PutQoZSS2tDAqOTwFHp4gIjb25we3i85W71eWsxmAXR
8EKMqHw71jNvvXC7dxkCDX6yAKTKIaHpCYh0YTEJHKJIjsGK6JJKMUWYroc69/Bn
LXLrtsGgoyxD7eqKJbojWuJpjit4Iiyj3oWo+ucyw5/8sjMJIcLuuxzun1mXhJ+g
HmnWdsZHbYkHNUDRtSnZrlsxeu2cP3wGlhT2j3BBF6qm6O/4lYxkLb5EPWeM/Dki
lglYwMvZv5bxJJOlwoAnMM/B+2RXzTI8eyyEfqERkzGduHmJEdm/XxMplIsDCuOW
KhH4dt8S3PS0PzMvpgNRSZNFSKyIVzrw1jHLAQuUraNmf+SR8n0tmoq3b/hhocD+
l/QF9S1pxfzW/wWvWyMf1jY9nt4YRAtn/UY26W2FMs4Nz/9/JHdH+iWJcIYDXnd9
KUjqlP+hHbpRlfdY1L1u6xV8PbNDV2ZRR5h3mg7Pi5FEAdzkD5/9kSQqBrsf1Bqy
7i/D0GWnK1Uw7B5ieYBWQ8OVU7Nu/h2PYu7cu6Q7HrHqQNnW26Yx0LhBo7Z6tOwj
FJ3LWWaKkNf1KF1seWisXjJ3ND64BrlAJckbrmtYLzdMRxAtmaIUhbidHly9wsi2
yNAbZe5NNRpK2xHmtJPQ6eacv1yXPsWbkVN/TBbFvYI0rgSV58ScArV0cxGk7RM9
1uS65J3iEK8SFs8E+gsNqpffps8DeBQTfKR18I+Sp84Rzs5WQLOrD/+shkO4QE+I
cTB8aMDEK2xzFoc9u4b1HsGVLLQMghfU0iPLPnTqBk7iJM8B+k/mDYxWMWFurbTT
L84dTp7dSt24jaTrwhEkHGu7JQ/sGBambvj4YFuFlWOJ73e9NiFkOC32F9En4P7x
fjH5LXDIs6Sr9t6isHlaWuVWWNXZZjFhp/2KcyfQxccrvA48gM1G35HEpTbzDeVm
gHmQYLxPWsflg5UNVLXnXmRYbycw/kC157PZQBI5l9RZWpUdwvRIFhtYDVLc8Rzn
Z2X1Z7rsZ96NEb0Aocm0y9eRaoqnHY376gXJC3evQT9eeUBLvEJ2P5hBWmXeNtXs
nPJDhv6YWn4s0WZ7yG72lOkezPkzBdFghn76EX7wzuEeHmagcGBNR8OzJhaKisRI
T1aFN6WIP9hZkHmRXHJEhHGNonx0elUEL4BzzNbrfpUfwDTvfW2m/UHKCnhff15d
xHucqcCqfxL+BI8KsgoWKk7zkn0MboSg8Cr815u2YX3U9kEzW7RSy8HVvnK1VtQ1
U4NdaBoivr6NmKt8fbsSbbm4SkgILn7e9bInX9QpJrEsu4k3+O5AqFbriKoA2MAb
AxEyaMRvr5ZFm8KgAEPbWaKC05KbrBvavbY5VCo1oBXTwtpiZ6O/aAMCMMmfJEAl
ZaOSQC3cpaExFs7IDpr8OmdhdXBomdd344sh26L03Vp8Esfhwi4hb/wOeoyqSFw5
mQsWDl/MEoAOTRIjl+ucMkvN+o2QEmOq1OeeWC+bYSwm4qsFJRxarvszDygpg5l8
9c5b7GpHEBwlNHEuhr+sPwaAZLpw2ANFMOfTgou6Kf5/EdNKFkgbHl1IQhQr78rz
nHkB9u+VZaTg6kvepiQT0xC62QwciwfHga8tU3wpRfg40plPVaH4y/Ma++Qeos+o
N6vSjXvxVu7Z3nmdzeS98a1evG6/Wqvdf00p9wZPTLHDulzY2Idmgm9RF5NoHBZf
YWXU2+MJ3TDZ+9le6XzAPxK6jFfbvBNuvT2wNipaACLcp6dejzY83lAcEdzktzv+
37ixs13oFn1QiViJDo4QqeHzAP7icugKXSwBWqh614gNixbh6aypsFkYospeEmVv
fTxDWgqx+J8sa1KsvdK9Xv84hZZoo9JvwLfJcap0kKHmv4M6ZjubOW66qT/+J91K
QHy/MXs6fIp3mhLwbxDC6Md/+OY6tmN7oCx+23Ev5CevArQ5yZtnSI5Mp8Bv5kc0
rYjD0AsZKHgzS0RXR56E0pgtMyZlkHTCkrIugQZPZJbsyNxsS64tmQDbqToYK1tX
Fjf3amc5H/Fuak3hQ2tYQOkQJCz/HG/0gY3cY9USv9sUQhZZ0BSW/aHoC2ONP2r9
k+RxHt8GUr5Lav3/GCYbMYmIH7iehevVt9H5Kq6eFk5qrFj9YDpV4HtMNHGphYPZ
BpQXxvJlYxZ/emLgHAEJSDIRZQjrDUNk4/n4YhVcwNi2amFathLrkqIoIIisq3gX
xZgUf0i7gSblQIdDvXqJuS0aE84o6Buuqp2OC/04VUAdHSDRt6jR59n53COGUdDa
vU/DRpcI6Vs1M65eNE9TuPrXtPm3aOtcpL6zSONj/xD0V65eWBY41vILNnVFBT2F
JkPpcrRG+5VKJquyf/8q6EkjddpaPcSaG81G2mtLJE8F08uOZzMfmSByw6jG9mpg
8RkR3E/ZNY8jMr8B2/fase6G0qq88ZJFzr0PoTGz21w9zF2rFIhNGpkWoAGcXfa3
5H91Rt1wvszAN6n6e1EQRNC8Xq4lOLwe8tHF0jdzzPivKPRBkQJNcdPjjYsUcogx
ZKlydi96P3KFZDCaKmn3US1iel5LUpscBLrIBUj2FHTweAdASn0PCVh6US4rCTfJ
OB6wsSO2mUDo3Dmn1Mba5qiw6Xtrq1fi1MWrPIjTJy0t3UdsY6TpXKOv32Y2b3HP
SaFPtpT8BitYxbowEDlq4tZBR1kfQQ8T6C3Z4hTQC11Wdovd2CeFadoxhogmlPGD
OZbSt+Ue7HNdQXr0ELlyydY7JqLuhZJE+YnFJxpJgsPhkC5PGmcW0n3RSGpZdXGz
OgXZBjV4ZK08HD+wJmxXPfHnHLarBMaHJDh5gCGLW1UMM1zGMQkBHWQpZ6Tq+lT2
kCA+2sOfp927YwJ4iNVXzgDDpmNYMOHu3ZRnHG33RFDzYkp0hdVrdjqJLzC385vV
4I3n3dOxBXpzb4sjNLYjH2Q9Sp5puzgc3qm4TdOESahuPb3otTtegrJQuLMqM2Vn
QDFJmGTFYd8185I83/7NVLLwZq7LiAD0iDaNWwPLAfPOSEV8yNAe/g1WaMraeqHy
FbtLgw516uRbsKqa57nGm7t7H1duJ5255ineCSFMsTtpvgJAFfTgRXGdXa0vB2jO
k35I8bbTUHgRko+KE+h/GN3oVT5VLweN9mpXHG+o9j5Tb8xwTsBCUfprJrxWcRB1
Ds9tY93S2FrDEk32UOquEs3z59xrQfdTLzXJXbqfMwr8S5yMhWbQwgVgGd8kEJAE
YFXtEkGDCHjC3f6AAZ977aDw3JbfPpSU1pMxV5FzibePLvdxmPf77KM6nUY15z/7
oxvoPTPGmlw6EXEgj03cQERWAVTTfTmwsaW2QAbk7xHFa2QPgcjnne27yt35mmlH
5udHM0X3l9zKjC00fOpj2cdHLZVLZOjYTpQ9opxSc0G7dW299dHE6qg+r8vrwUgK
jx2a/g0y0qFZD6OHDxuE8fYVeZ6wrkXJAh/gW3Zm9JH7uligpLHmLGdRW5pjt4PA
e88eAmvBMD/rESwDKYuvja49N0nZ3TXOft+lC2x9CXg3Waoi6fC/GKMworRmwlMg
qvb+aEvON8L3h94r9NcnkfJ2cerHzgZU5SvPACByOaaq+DFRcTkUtn/5238v/kty
/XyfdLXrcIMY5/cVzynLuio0EDZccGjmEemZYR4wm2a9+Fp7X9AdXhOXnO+/B2OR
clJwuUFK9yj56SnHq1Q4l361lpLkevvO+C9rggEikxt5eoETdLlYuExYq2aqS9BM
sd2RTsb6DttdtAuZ8WqBGQ/gdG9sP7raVUTNNoEtxNiWd83NRaoOQWTwKR0nRyJf
2o9eNE1gmCjlTiKw4SZFjocp5x0pCEowRO1CxEjpEQWohYNxYNuw88hDQGPjJYH9
KSC61kFLCjNO+SPzSeHPA/bkve/ShEzJDvPGW6EXaIl50YSNOq+NbSOe9eU+tAzN
2RJ8tis8pRvifQYbECq+yMAJm23ZLgNKTMIg68kFfGYJmqqWzceDYHyVgYAgCmIS
eI75g2cspge2pYNhnTOKwoZZFI3TLL8SJ9N+PEZj+WKZNVdkNBy610plXZS6WSp2
DAcypFy4YLOuzEfHmpPOF3+a31D8lgzsq3qmF51b3b2Hh9krLGUAxgOs2FM8qDsy
yJsDfxruQTi6xuKsD/cWytkTasAZ/OCASd53sP+2a2t1NCHxx8+Ye+mYIfHDYC66
JG+d0SZzVc5K5N3hshNkCn2kIvpYdZYMD/bEJvLsf3hFHtSbTB1BQdZ+BNGEsnZw
DXSBcS3aroluvQiHta4RZlH2NwLBVpehbXpoL6tWF36KuPbYHLh9rleP7MPR6oNI
k+tZwyUjOcXbRH4PUKtJTcvLxnLySlxLAffbMaqErvO92nlZGH9YgcLykFtzDpIw
JOKEKHYXffSoxn+9f/a/ooqhyhR3Ex6xSSXDhnFm6nIGvl41qrMiE3tqlalhPjba
Z8wCizO13e/7fVpxOrYeeqnnHJbzFUhqwnryhgUOBmSiTg9gPDdrVquygWRHcGSw
v7ee7A61IIC0cbb+mcMnNUO2qT2C2G5e27h/1qxAMBli3DkTcLCYHtFJm5eIZcg/
LUfWl1m9DBYMDv1Nxvc7G6kLm7FiN+jd8T8PFdn7+uRFiTQp0QfdMsiVNQUHtOmM
wkIQgPrUbon7p+tvWMA0abKEQgYuBC2t/vtDENmY+gxd18nMTwkszTVJ6phI9hSC
3L2phxrh8w8+Mx23Kty9oOJaZqT5YjrEWkJDALTVCXgoKeD76wUw3qqI3MoshIg2
jtNZdHUm+r7Gwv0i7sJEuJNHU+NmSFzluSogugRFnVYGDTELPlUoP6Q2hlbsrFkm
ABYITqdg74z7gl+BaFNVo5fgontpy+mJ7TShnTvxkErCyJktaJ8+ws+UDKrA+DS+
qyfZAv5TwDlq3vZ+fmYMHrrmqUGxutqU6JHmlmZ7iTv2Ta/p5YXw180/rlzj8EBa
z2ldE47vimgdGcziKIbWowvyb1B0sO3U0x/J2JAPY4Vn0Uvm8FXIQcz6d8gk4Nqb
QdXvk+u0kxMCX1yek2UigAIW1Y/GZ6s6JJDIsVn7GMeQGFyuFtaUPh7EBIixmGJw
2fm7siQ7Bq/PB6MfzALXweaexJZLfrRA1Avj46Y2H/Bo9IVy2233tvarT8eiouKG
EE8FSbNA6FBkxK3BZ2599dJ3rzn4NVpf5w8mcHqfrM9ykBUNIQIOi6VXBz2uZGTa
19V+uD5v2m4luGqucRJzNFO66wSczyeC7s3LUk40C88lxXgeu1Ie2kaZxTFv6Dyr
OYip4DTJHOG+V2WjRMF7YjTVWubU5RcsNUwzZ84sIP4CNoODIHC6E8gDiKr/XQ15
ojnk2UIh6qahwUJP5zX9O5n2FCkIO/YEw+wNQLGfS5caRMr+6hBYZhFAZ2hVXSXK
oi6ptLaCyhSpVLyeDtJ6yYI8hhgNi9++3czr440sHJ8HvyloEF8BtP+ID2H4CXuR
T6j//D2jiiR0qucYFYdYXIOqcWjsFsCsJSQpjAXI2mgoAs6tbkLloI6hPieEKUMB
dm87TaadbtQQ2IqyYw8NE9p97D2H7srrh3W5k0k5ntSmDib0hY/dmqGBYJ1J4tZ8
1WO/rx6Mf96iHBndOTgS+8puWTwhw7T2hsMVkjkkBN99Bnd9LGwXlvj8k4uX3VNw
6CITWKC++PlvJwSi8yMq4o7FIC/1oTQCXw7hv/QtXjc9MCSi8DGB/1xJgcdCPEn8
Ig7+EvfE4G/XbgkJRXL1iml3GEezJNn31scsTAYWmlxEz6UnPxJkw/Oh1K2mB3gV
fTqWwDv7WdhBn6y71FBBt/jCl5KGAAU12OheL8gTX4/Lmrq7UiMnoCo9OEOmhCyF
GM2kLCWpS3p8d/N0MRRfgFCQfRUi6vYYEvDwtXrhkjfVE1smSkviAoKOpCWCueGf
fettYnXCBYI7dBc27kYQtCXJ2E9W2oKnF7X1TXEnZ3fLw445RSBlFNEP8ETibVzg
IbyRrUtmxwwo7OSJzCicOBhU29+8AQWyYHVxvQy7arju/++xgSymDz5FnAVpkGze
D7FFGPG7WNwk0CyAkY9fqu1wOMdz+KaLKTfa6usEujOhO0sIoqITbIwMkJQr8gNN
TBRD7104N45opSKXcxehJq16kmMHP9apb6LoLVl3kOafZTF65CSOSpy6LvOySby3
3y22XBQXoZXKJ1vYFEEFlamL+OKzsPXu2RuVUJJw6tF6GoWFO2/312l9JUs+sw18
cjQLJq+k/DizJGiVbh6YiCEfgkdSJyfquNFKPAb3lNwzx0sqGXC98kqtD9ZflqrR
e2ycfwQ8ns0UQZneTPLvbujbF79iwWYypJhPd8vkHnPyb3QNjc2C+jvlrmi5QS2k
KO89jhemhJqQZ5a5MQyQYjp7M2dgCfqxrDEESOpdFS83OYuKSTkkGjzww9Ls7ig0
eAsWrrz1FtXDSnL2/i7UHEmG5/k0wnuw+++30D5JWhBU7s7MkA4mVBr6aCYxVlGu
zKxPB+4kL3sB1eR+dmx7CBcllKYRQKZYIoGTkTMABo3WEnb2lnemzD3fJvwPB/z7
sKXfo2TyBBq6dKN3ofhiGRVKY8WuLV0FJhV7hExYdkMWsT76GRYZhgzLaO+n9mZ5
b+XnCgKyINLDOYH39LxWhdnu762YOgxHD5VZbTcJQWOhjdMNT2FDMTQLWRVhpyc4
6UDUa+JbqgvATOEBMjUNLNkFDlF6V/1oh6ybJl3YK+mcgRzs9Gg4c3NoZVlI+O2Y
VVmVKYsjltUYza2Ir4Eo+EaeLcj2pcSKNCibOt3QGivC6kz/Mk3XZUu/DYtQyond
tmvwfDh/msbgZ1GQjOk4VVNJlHj2asOz1jl+4BIoK7seg+7/tLnn2na+Dqid4f48
Uayn+ttQiZo8HBphaRGOvRYGDAissbgh1aIzztkt2161Sz0HfPUQ3K5XOe2FbBff
dNLPhYxoBh1KVGpJFZm+FTGF08LIl4tX18Jcan7QZfJ9jyCbC+pE5sq5imgO2rJd
TBYBrtHkP7vmtLuMLc8HDWusdx5/jVh2SoR4U+KdJtsM0YAfxcW1kQVFJmSBQFyw
Qy7Mnpt4It4Y8ljGbgV0zB1z11gHkMZRvDSFeFpy6J06mV+/IXZUB//6rTKVW1BO
9Iv+sWdiyfXl8809aNAb/bAMWV3G1My1m97Wut6/42FkoElMtoGK8UtUhQ7urSya
XPSFtUMhy+ddo9v5etj2i13+5nfUuLFHAToxy9fbF5AboG7qyroCXTOLUTFkWbO6
f+R/VgVEfduem773TUStItjFGTBAxBik9tuROd+whwbkH/88HSSlNDt4WQ3DFFll
Qld2avyITQ6+MvqSRih552n1dROcjZl3u/eLiRctlHyz6w9UbV2iWts03vHy2k/7
85Y97UAQ9N1GNCVAfnx5FO7qa7Np34wVoyMOUiJdrJrIoijOAIi8iyUcWe1ifBwM
aanrF050oRvKtEfuhznVJDTuD9I5C+B7ziquPuZo4OgixIYFSkEZWUgEalUzxqMZ
rgeRY15jLdoFb7WYiK3ZilIaaMQq08oZchi7KPEklI+fou372RoU28OQ6619g/o6
5Tmv0032fFXeq5TOUFDsxZ4MBqmJtCluYvAJ0mlt+JnSo4qeMKBsnuvn44y3YWpc
6RJoChJ4EO2y9lF05lad/6+wzvF6B7bqRdovk9qKmvvqzScDCJmy7QlJgoBBbdB8
gVHjHcgjEjqQV7PZLrUXrvynX/3dEBd+Yl04plvcF1pG7pMKASs9I9SFDYOIZU73
dUPGRE4ZMvWR+XIesWk+zoa286ctBNDryPSk8/+bXt/f/Q7eIlwG0FRrkKba4uHR
kMyFUceeqOSAHeZMDgrOS3zfuo/iwtBIBgTmvYjJ9E+dqbOchpimA7lgjs/2M39t
3CAIF8YCK3j8TqlHIKnDNeJJoA2m8xwg1wvhxCqY+G9tgPvNfaxHiXEqn0Ss8jzj
v87sYiOyczXalMNWPCJPHEVbbncl2aDZr2/a+BVXxVMGvDn/p8sn3X/gqFtSPQAS
aIsDSnkFZz+H/+8pwY6Hkm677xhejc6x2qnlC8rMwL5qO5yo8VCMQWTb+6f0SdlZ
gLA+YBcGTtjWikGKjIrAC/aL/jJI8sbENg0k3VKj3YqHtWxxG01ZL34sbsvYzNf/
CCQHV/oz0MqacCsMhC5YDFQRtXQ0duDwTVd7qeZP1ncDsttwrvLkeHPtdOEog8Vk
+A2hi6yplvKUWxvMOsBuDaDDjjIQYRYfuzgMt3u7zqJqu6a8JX9Hf8tgVsUW1C6Z
H5lypkEvpzFOEIif+xOWg7Nli8wLTgZqLcRgaCSnhLUEvsaSLVC7bBkF5blJNo73
x2ZG9ooleE8E32VJgGsYI/ggQNbc+o3XmrHp1HtcTXUg9H+/wUDLqmidf6A3xHO7
zNrqvj2gycoPP6agRcsE0Uy5N3Wf/CLqa3VeeExMu6sE0tmu0VvhpeiVpXONoGzu
iOvqc+rvPBkoWJuZcmJHGyu4UcVFo2yClPA0YnVHNju7ZBfAGrko9p7z4j9q4/0L
dujAD0uJ9HYJ7sUWN0djet83Xgn9H38x3bMaou3dzNHbNULyH122FBNegt1VrPcK
Sn4jp87lvumzXBv2Md6e0/XPSSZdm4wBZ58JG0zNBADZpZB5GRLoJ7vbeEIG5KXb
HnWMysNmoU82m+fkVFy986OhXD+f/6oIyLK8Tn4/70PGz8y82NwW3IQ9WcQQHPGJ
6NMQm4iuRlytGA15qSUV/fwZIVIXvI6RcocVUSH6uySfli2KEAQ/9BP/Yt5ZSWu3
UC6S6GhmKrONm/XKAxhmsjEQiLnx/MCnn5Xmc4RqvajKQhXOaYG/GKTUJ4d59DbO
4ArbDj2QkbjsNt9UQzteQJtcmSdnHNLcig4KbQk9GwUzjlI6noJIoZgJDXO7YtKM
tTMafw1OFWSq4aUEBUjL6B7gftWtX7hvsKsRoOwlffaZBjqK2Fxpje2GUI9rSv+W
JE6UrKSv+9/Y0WRruZBWPFHYeGrrPeImezkgXoS31/tL4bruLwoG9ETWIwfsNWyd
vULSNZnAb0Kws1NDWhrhWrqOQi/E7tgUIibaraI7WfU6eK1XVYiVBngzlHmqJ4jU
fOf3XW7eSXs7LSv35OmMGLJdFpfjxZiDsgBjXcSUgZPsZST5jw813E77/TpPM+Mq
Uaz/uwdJ5sZKFnEXN9XPE0sYhWmJkRrQnCg/x7Zfn982xacnI3+Dc52cLJs9Umpw
iu57Qbey58ha6eSWZV3wBAjwd7P+Q6IVmPzbzlsYH36o5IWbE3wapFgaU0rAyLeR
gdnSB+U3MQnyI0hiLJk5QQ+evi4vo/D5T71+6u5EiY0zeK5SxwcapKM+CRczD3hU
jS1KqVRN+tsxqbw/sWQoOl7tcl01XivwsE2yxH9DCru/Ud9aoaaq091wuDpuintM
B1WBJlvTv9tHiXXFYrWCu0W9WmbDeGw+Jb+31WiVIpw/YC3ah5iVXjDETiLOKYgq
up74P99cAJYBjaqT9xlSsS+/FuGi3eyQO52CCcHFRVSpi+4h/Jqpi3IUvnBnyCjb
0kQM6hTilSe3/+r9dwCT2lPJU/Vil1gLCTCtWY0YPzDUuhPUVZy2ZnwhY78zajbN
dFdqhKcqRbGm0iM9PsogMLUCc57L79yZa/2TNFks3A5oy/xco1e8lDO8aKM00d1j
wfxZ4zV1yp0+y5zB9IYavzeM1jFpUOI0Oo91tsmLYb/887ARtnv2NF6gMlmDQNQW
zR2ZTUPDkp1dJDLstwto9rew10Fki7Ir7tgNItSySa7rWZLmChQzoF90p9w4KepF
wtZToBXIMxDsTO1AC0iqfRhBMshQAXjO6QTtAyD7vIsgzEC470LiW55zOjrON6i2
ZL0pxJz0L9UltH5u/prbtflpCZKA2g1lNIMpcCCq9zxU/VfiZBq/SjizyGiiPUUx
OMT0xRC8X1nzTWAjIXQPOFTNVJNl97LyOGkUy3dM1HxSBzCAi1PrYSfGRZ32JFDv
PBfURhpRWqaimlJMjIgfdTezzgA8DIv0XCFwc671ekQoUmSPl+SpvVP1D27xtOO/
TvADjeAnqBEsN4inkaKV48EEes83tgx3gT47FwFRxOmzUaY+tckbXhrPVhaXQtlV
FAwTbkD022VrRw4rF0MDFC5LcPuyBgxuC6u5AghxdvPQW+iNRRx1hFDWMqrf/mDv
r9+R4BlxWtaMFDj+LFRW7fk2fwuRlzmk+jfqKOeDDxpepPyXd6fWo4G8rmX1cCPF
MiDQXy/7FAkEMsL/Q7Pp0Qvdqqo2UD9EmKIhL5EZCq1SJKltUPVrrv0N/73mW1cJ
pzoNp0LaHnFoFCyRRu+XRuzKjMI1L0hF9PfLXYOwcxSioFd62rh+lzEZqcWSzHbb
cHYGTnbm/C8a1jPVX/I8RFEmlsvHiXc681MM9II/RkBelqMOs2mIG8/a5c2Jk0D+
OuKgJKz1gA4ine/6a7fDH58Q0juCSXzAqC4nZTvHUYl06EfW9c+24nSxAIC1aUi+
HSXO+PJkoHkEFd2k33W1lg9aKSR57nWJc9himJdIqB43+KYuFzljQiUsRLjaMio9
KPJ0rM7eRaB8frULn7dl8G/8gQuOlx+oCVuqpldr2WOSJTUpQ5mNOgwDH1XaTCyz
+yeyzHQowo/JrS/kt6O6ScJJ6+OK1+ppac3AQcLP5Q5/+PZeNuyKhqWtWFM91SoK
Zr0vk7UUNiEWjj5/TVeJ+zBJIIgd2mlzQRYoxaqn5TOIUAAhFZGqboPNLdxgbC4I
F9Iljn7yAOtdwV4QMd7pm1X7hSIHgHBwFTS+GeO4Eh3uwJKPqruoumMQQnG06WpT
r4Jvae7Js5GKt1fE6vDxce6LLHngdoZpTd0TLqFYRaQeawG9wizf1GMzaX6boixi
FvZ2ip5BjwPSN0toK/hi+FXGrQp+vFW+923yF7vHGtq+t84OCpBNlwI/ApsUp3+q
8k+RlBMqznYbuoNmafDMlLFE0A3f9weBSMJS8iz4HtJrEI0LnJtV+RPEkT4+z9Hg
VxPe195pdfVg/Hzw3BsHMj5lKUnabArxT5Ap9+7CSsXVEseV+xVo9FY60hyQWGQA
4OcOUiPGvmuJOcE4xG0bvXGUUBNHmTwaY4rKW1aKcakhIfRaMY3Pj/DHdOqHY5oy
Tt3a15zGLCIMo3sZb+288lGICXZ5PJuiZjzg+m4lPQNvECd2ZeGJ6zTENj5TGa9X
7s8+QNGKH4+hwJe4H/Pfhl+rbQNB2IfvRRmhA0V/9WxXbLFbfUSmIAKqCtKOfuIh
lMKnk69cJjtal50h7mZ/n7ZCryCo+l6nH2HUy3F22oqI04TXAGRqdQopXxT/vC8Z
hXcIwf1uwRQxptGfqa6iL+YZUhm+SeevcAsJfUScrLYcwewtdDtindfpFvoB0wGx
00XYLsEQccotIquD/IbMOmCcIuEDJ2PajLyGPPvVJppL5eJdabj+w5Jhts5VaQLf
yqCGFgbQshguuHhcy0cklhuP3w/D9YTd5vDOwENlbEab1UsFY6WCj2UESY+N+GTH
vVPQN+x9lrPb2DXY9VI+F/DtAMVisAoJrjHArqAGXCiNfMAZHm7SD6mT8QZTawu7
bd/sorFZsKtuWsfqO2R+UYsGIYsgWszFc8icyumb0qZNOKHavpy3RQ4NalvnF04S
ihHOqRpXAGOEOxP16xAt6xPf3cCSG7+dxBBAtZ5tAoTqLMi4KeH/olzRRKbQiIct
Icmw2fbrTOznJvsZh16UmGD/9euXvb4XLBBWW69aAuLd2dh9f3xiQZX7NgqnDjc0
ZeeiJ6QK1aynBNOPZe1CjawVRd4UE7E319NqZFBFlWTRESAbGGXaaw7/6U5bVGG7
w3PYwMHsO+NhNt1u8ZShBOrgDy9VsN2ot8MFme1wI2A7DWmMOmzsddjFjCRBMGzi
wiK5rSJgSI3OIG2Oqwki/ou7FTl9jAQHCLXRTncyNgsqFWLeh6+YHVAAslTs/p9J
FYs1S9sC6MbOEEXFWP9KBBhOZrantQ4pltJjdLh0LR5KPkoPqCOCeylWhpqB06HP
Z35aiglolwQA7/w2vDj7T1MXEgBywby2wEdDJqGGk6DZ3kKu/jPU4pdU/f+/bMRf
2DHmIF3VRzCz90usVTUOvHCTBELJxBSt9rOvyV6zfd1+34pODTveP0fJLz6ZMNoN
YctqCCvPM0ncFQO1+cKGLYpOrIOz2H+kZLbz76hHNemtKudcG4mgB2Kn0yvyurLl
/T5GcB9ihFNoaTmDCRw6ZtfMXRRYr+IzYgr2R8iGIjSpBE686a9PvJCwutLjMwqO
TblLB03LZ00VctHewLN+qm90aCSUFSZve2pWvPoFE91EvEzs9Qdkh8Jr2WnPy7zM
+J+PZobKCzQxp79s64S6GNWAjRmNzhLwkgYJeVNV15q1D5tYn6AddL9qMhCvbCW3
CsIFWUfgqn817ET3b1wUMs9edX74lMnc9fslnn17FVaVDU8wtFV9Q/t9FOwL2DSD
xuUHhOURXjCvLHTt21Spbg1fQ5GSrZpXjPgDEgSliPWP15QZoibc8ufdoPM6UBDg
3UFZznpF+fWbDr7usDMlxtnQKGiWxrSVhSZzSxaVlVY5NRwzuhhvSdK3qSxX5iYI
0NAvioeYmAQLy3IxsbE8HKXjAIaEs0RqZ8ddzFBGAhOc7+f5Ou5BEn5O4joqZbAM
t77bkNQbyZ+WZHVma81nTmxQHVEWa+KLLd/2kpQajkO5HW3Dvh3q/JivWkhfl8y1
Sq9KHlQgdHWgWIBvzSUmVh5XvijGMGSDpI/vnml6I00Gbx4qX5G4kzLVuDrC7tqA
pkXXJambqWn0ioDwR9BmknBYziqBHqP80qS4tJlIRdj8hf2jao8GlUG6ytyjtSNZ
s38kMY6+GFzVqgrhj+LscYFxM4e6nPMwIZg2HyXoO+AobTxZF5HO+DrCaUEvENTf
ve/sumCT5pUCUlrce283ZWUnDzve183k3T4oo/YtNOxJtjrpZ/WFvcbW4fFH4NvJ
jHEYwS9gx0UGwHLGt+bF7TVVMg9YmMUfSIrA56Fp7kg+Vt0Wm1QRCsE1roWHJUH8
+9CL3pLrkDRlR9icXEs2Q6GxMYFfuwWDT4bDjH0uYEgv0GuGc5Ql8j1XUhyk8pGA
tbAHdpqcGb41VCuaYhhOv775VdGoV5+ozCVnq0gnmChkYkbCFjUUjAwXm3Y3nAby
ll7LUjFpCF1lYScKccvTSLjsjjpHjJ2TX+B/mnkhj4sdlOd0iUULPmnuoY1pnxVb
2s8PIVA300tTrfFFT0i1pe9I9Eelk2Crd8C/KYt83JnFsnlr7ZQkf1e8OO/Y11Kw
mvbyfvUz8d8QU9SLRxJko2wWebc+XNUeyeTiyqW3sh/rJS2E+ry79SuZRoQCOQoX
tnTvN/mWGjyGh3BB14oR297RAxXAHPkGoiv5rGG2oDpn3wRBqAn6hQU5s4ghkMOJ
oF6+SLp2bFN7td4BdrS0YBzt5AhLQhOLxv5usMg783R4BCu5J8GzWaXHX4PoGcxQ
QUbCuiH97itzbfUMqrf31p+ou1R6kMvvWGlaN1ojoBWhYr5pGKt8mD6xZDmZ/+wq
wlTpEWO3op8gdf7DIChY6xgOqpks5em+9n6y3ttwJhdX0SZrtOa8goM/RaxKiXX9
JHr3j0iropK8k210eeW2xKbG5DoTODB8mBYNCPpsKo+xAxNNxm5qO/R4dNVGnqjT
pQ1kHEba5a29xbTCdWD+zJssr0SYd2ISygr5/an04ZBD5dw0pmm/NoJZFUA/1L7Q
fOyT64zjK38nP6sR/UmjM44NWb2FIPBFxhd7HBHJ98+W6k724I7gZ0MsweeM6Bye
MXYLzKELquVeZjmPNJLmiBJHiqZoKIzSM1zVzcGMY/kdmGVEtpkYKtpXMv9ixU/k
yLDYde5sdkEtTRXFM4MSkxpCG+hnxCn/OG5yRj61atZ1xFK1Ci6g8CEw6FxPUTcW
+WAQnkfJUl7gIMzNuiYhbzfJbSzv3Kj7HBGBpP5Ft9xAVIpsUoBWc/XWVOXYCJES
gXOhL94g1LcCXkqLVTuIewPRDZ1NSEhzD8DxDVfkPObGTNs6fWRmKHqVBZFLgn+h
L4a6NkyCzwxKfAXD7qkJyfVYH7808k2CwQUM3mAMYS87KUmYk8riC869318IUXMS
6PQuXDOofBO9Iu16sAMuW/m2t1iZ0Jy1c9K6+V/1AM7s9eZSd9oMLHTlhJeLPMva
8Q3+F3cnO75vRSgSJPH2TTykNCUvHR3MtNRZMMB++ZFc/upC+XBTSWBA0QJobE9k
OI3+b42/kBdOjRv8hHcHh+938B+23WoJ0LBKj7lq8Y2ayBxcAvazGz1D3oGjcamD
5Gnw45oNoVzHCCNM+nm3YIBBgPxrx7386AHY7sbAlbq03YyXdr3k6MsZNoOWflFq
SjVBKtwPKoq9DTwrbF4YrogU1v5Mm065/rG7wzAldM3M47mNuoPapaPP4z4LWpHK
A7du2gJgY6WaliukRthR+KVZqWQZ0aIMMD3yRQnWwTy8BJVJIyJWXO+qsdiFesTb
CtCAtEZDTBQR7DJ/vFyhGtC+fiSXZISNEtFEIiU949PeP2xd/ZE7wG/Mqo+dpKrM
nLL0I81ixi8GU+8bph1pwj8MsmXlCmKgMYInLdoWmIdND8X/HKKy4V0rtLubLCrl
QThl+PhVYXDXhnjLtFnNMLDG3lllE0FtHnD5CpiTjH6bwousfuGDAkT32wy+OMmF
d0Tcp43eJFWji2R6jGQScVc6I5gGt0VM3nkJIo3p9KbF8ESEwN+4Jq200NeVHBS4
8+9dFElwPx/I5CJHzMQXQiiymKQdZilMyLF0OTUeAuY8edL+w37+O8OuoWVE4vRR
rUyYaXmrDtVj0M+3xG7lLk4UJSDDfYvJIwm/jFuLV0QF/dfXBkPFwqgSCIxJ2zhy
xyetnwZiry5ZN6muxOda7gbXr4Ta+pW7BW9sZ5+O/cz1mGB+o20UPuHRtRqOQc04
MBEWDXnZvNWBDUZh6cBC20f1EYW++oq2DTw3lLuO91CuPyPoGx1X4ZTrZR4hvLl6
GOu5rvbJq/QY6QFLd9wQU/16JHGT5dKZjXY6lVXqyXPmhMiGK5ICG/wUaeua0G9s
3JNppIx+/69Zu2Fyip1GUL9YER85ocrYljv60BuHQ8Ttxi5xLOYFcrwQtx7RVXEz
fr327k3SU3rkv/EdPgj492Clrfkk/2B1lc09A5BoyujMBhqylwJFteDbANykv5cx
pL7BPs3YpLz3zRCGjUkCxQL10lUt+oWYpkBTqCbOgzUwEKdVa38/xsNKDJ0z/8rF
esKIw1QVdVNLGVsGZF2zdA75n9JaGCu0pk5JaKJ/F10ydM9WgnqU5kYM4fyGJmyY
fBz+oZfAAgFejsjMmA8aj9jZBRCGl1o2VM0GsmmcSRy1W/AdhkrkFwGG3KKkiS+U
KPnUKV/mfxIClInzF6bPSX8o9QPH/GvJw/d8Gdzt3sa+I0NKjjw6hkedX0dJwEzY
64dFix/j93b1Mu8Bfd4uKhJeerQaTtfdBw5F+NQwJZkl5WdYYzh71T/V8bUgmVp6
1kvGUhcNkN/oEeKEI5aMdDRqPsae04z8ctRagp70hLoN1ZzAcPJ0/P4xyESdRY1I
XSK2xMd3SOBVZO6HbuGK+JvzPUoI9bst1WuqijzrvhmCOpkQsjUxFt7WidnFDKS+
6yNk20TBQB/UkMvoqiMEiUmQQRUve26uo00U4Ylj060VKskeMLHMYgK7nlSQ9ZC8
PUv8urB8uPEJ0aF+Qgh3pAlLx/+WaMfJJmeNE95Epm1jAIO/L8HahFQ3z42X+Ikf
RUronbrsvPaEBqg8TNDsGxb0CwlyxCQiAgxFDS+ZDeNni4hGx6xEARghf9duxYMn
yuDlT0IoeVSrY0xgfR7BFsct3dgEio/1yUdWVdgaJQr14TAI4K8jgQ5J9rHCzlOa
h1q45eX0rauUTdRUPqAm23V2JpLCm9sCeZeGT0UgvzqDQdkAm/gRUX+xh1+hKZdP
JXK7j8wuSmo3QzNP5IvcyzxuyrN5SxDGLGCatohSXEKD23x9xw5Bvjh6q5i1cq5I
nJ+pvltqUdVMB1kjWtmVUzqD2jy0rmuHOiuHEnJxMf8fyMInRYWxuBPzcXvJhRJA
7TqUVSoniGRKvbNojUuAM+LYwNTkIMjD1qH6ikWoQW85OVRnA/d+HWYUt1dDJpHG
ST9I7fACVuUSR+EwPhAssA5g+rDfetS8Wvyr3wLMJBJB01WD229hMRK5wZ1TyNaZ
Z8q+kkJLf6MH5/A+TJS3te4tw8tQEwMrzNJL5WvordHsdzi+bmZclUcMoRE3MbOa
l3iX30epgCX8/LzysSuANRXtSpgj4b0hG3IYPFh3eTs0bnVtemfGFDPw9qYk/O4l
usGIiPF/65LTkjnk5+nOBXKk7TWVGBDyhey5hnocrhS/FqoD5JeWEukJYkJKazeG
Nx+ZktfAvo8AK5RqczNiK45c/KZb3f8MWyMa7VTCaB4gyobZleD/neO+tcW3+iue
+lAH/ebfRTXYaUSMo6U59Kv3ZfEh/9B8aMEDRFt7GRZZqe+zIqpAy7EDm+0oBfXg
v1Ldm7h6JFcD4tCTvi1Tghph82dLqJDky0UViwkV9e3hX1vjlwodB7bP+lGr5Ifv
/D8WTuv3L2Y/sOOjapACP3lQ1m+gtwS9E5Z4S1NQKWDuLkHuUWaiBgqWsT6Jdevr
xDnqr6CVwn+3rkoaAa4yRmyEU01M6EfppsgtuyE9HltDzsdf2KVahTzkxZkAPVCK
Uz6bh7/Ta4N58EPVLIRajI7mOTscfvIpYorNwXEBwfrxT06o4nTTn4r0Bi6+qMXm
WiNgZEIMDKSOQbx8dWsASluMQI2IiCzOZ4Vo7Dlq1kgJIo5Gn2SEFWAfYVNWZWWj
WMcp5n7+3vScKZtbWKWch+K8CY6VCnOrgx5tC/xdRH3RbbndwAZ6LHIENIWVcGZO
1A0dcfv8HMh+p20wXBJ77+TU1m8AHZIbmwiS1x/uTXOXUphXZRnFibPVcBI9r9xK
J3/364HiJBq7oZtEYnk1FADLjo3TnPASYScjmVzShanEqSoTJKSk92EEzKQyejL9
j++foF9R2v8yzxX9wft47VWN8m/NZK5j2p0D/vV0ZFlqLRBrvwrnn18hLG3ncQM3
LSNDqJWdbH7knzY7m7U3uf3eskqqlP8IwnpbuuBcU012XOcGdia4kEzke6ap3iaf
Lf5y5JfP1iAqMA4xWudWflei9I23ziIjDWpwdgTmXs7etT/iwOdFyoJBTxz9/KjH
CxlwJ9HmZYgdzvLPYrynMuqN9JCa0an51Ps5+wkQrbVGYIcXY+wW5MWmWPArikps
bdP1XFXntqXHacwOmQ5t/CIV0sHW/kgUjJALvRK84s9fvdE6r/ERlpDtzrMT6Dm8
fKpuRpVlO7xezX0+qTimrLzHgxp/2tnJZqirGu/3K45apWU2G4ECaVO1XSh/khCV
XzJ43EP6llV5r3syBWNY2PDii6/WsKAMcinWAHRW04Oxj9MkNGIMbuvdz/B0VAvK
li5HQM6izaoymSlHJ2V9x+lqYZFlu+Yco/WzA4xvLihl7q+Yci/9pGeZj0iKrzMf
2o6kV/ucywo5SWBCjQG2OgfTPyaooxiEUyWRL+v0NbSaxUh6VK46gSJCbkDpVEYL
xxaosyD9ZsJaPqdQvzf7384tFqj1SKySnFaPhnEZRl0cgS6SSssjYWiR6s7d0feZ
Ri+JbsNGWXHNcSs81AtiTVpxRodZxkqtOqPP317VEhhzHGwPhVZeoDmzQV1MEMeZ
zNRA3vin1XiCIPrDt8ccb1P1QDMdJcrUxVQLald3WYbt/+Vp+2IZ19S+u7hQkeAc
hFZsnKeve8oGpbsoWDayBCWb2oiUuQEkPgY17szoB9XARTd92HzjKZT1xVUbG7oi
rrRuMn9hPJtSlU8vGswzq6agN/OUIu7lTRnTDBCczqfinZGnEGhvqLO/aS7PZz8T
SM+/5WsTMwU1hBh21vpjVQE9QglVbJUmws0D8WfSCb5gtosxq8CM2wXohRLzWdPG
ANSlS+UTL5B7M4p3sjZ4THg9b4zQZzWzwINd+0LYhDyCnEGSqBLoGU+7JxLIMWYr
tOgDXwk6kYig96DQ5HF+ZQL/K6paGJv8PWBWDxHA2LY9jpRkFLLg4Vae03a6aNjl
g+9+p2bkrVJ5b/AnCXVhJdI6wWbzgagnfHF46mAeouYThayuyLoNo1sVP4iGOvRS
chzKYAX+i22NvyXZfMwAMLjrn6y+Z7xZOEyUqTXx2+yGbeMa5u/D4svL16eruf9e
Y46Sfm4htYBMAS864gMv65HvvXsWhMlqIazsy9Rjx+ExSwJSqKHjHlYaodaACABM
zIV3VsH2TB7FgqcP6SGslCdj3HypSpfsHRqM0VsGAMWWPxFn8jsaGxGet+SB5YSW
1F7cXHOLB9STOsM/o5G+4fu87gXBWuL3kZRdVLENCsQWdVbAb2ouNoyFSavCL86A
IG4NuvTkw3kASoYb0pPS3anaxL08YGwxM56GgStEQ3l+jv/M8x7ByGnu5cgJyxk1
MCqAUuvhDXbR6L8V7RWL1i8uYJBKD7ecVg4aLV+677xHFGwChvfBoQbhHxjLQkzo
NanuvSMlVFi4HqkX30JRMMN/IMPKzm3r/vRXi+U/qJNHxm4z2ixslscL+4utElad
/JALg2B1A5IZpRB6LfCsgYekB/iXmAkBe56SX/gPSaTFXEIoEirogdx0e3YlVJhy
dHTSJ91v8kSzw8pte5Zi9E9KbhDky7Ghx74GFQwPUPsdsH73u3ItLG0limV8ymVg
pIyw5yqrO2q5cUgibyfcq8FVBcvjSgO/O7eAYem1w5vIZmWIcN1NeM0tvpRgLz+2
eN6P81LR2/t0su53JfpuyxzlV8sp3HvG24w+cAAoR8IflHy8HPzL75g4FB6LHTpt
Qjlqf+NWfuxvD/nYaZuSuSZyJJgXzm196ipDzQ8rSA/vmnYv+rvjNVcaQbPWJ1f8
1ODnRbLUWrf+8MaQO6xW9dipq4uL8zs3pIRpDnf35ccNwutTysuLRfNilrWIp/Qx
avKBFOzReVStvkUdjxpTdJQtJGRw3l6BaZOzPHL73pkdcxKzxS/DTQEX2o24444Q
nfFjkBGapDxeJlQnWNPW203oiiGYCii519EHcbkR5DI/qvn7QpQkVS5Mvo0Y62q0
WNdvy2J3EvEnx8rRW772y+EF5/N540rE2+WO62OaYAiq8/QDKdNynS4iwUpjkFwg
vFz2bMikSulWaEjPtxbg8Uecd1kki1NngNGbqigC21/6vg3cALQ1ZCL+0s0z6oiN
v+AMcd6UOMJa+ni3EUp9+gAHYVJ1hSmZBT9uFDsKlMpLzVa1KvJv0wSM1B2svXDh
paQ2kbjxlw2l1/Xzl+Xn8ukuon3KZRDDGToA4VNbdBZbHb2qYF2eOG2cd86d/KVX
25HOBf9zYhM39Y7q0B1ArugNaVYOV6pewAYz+1Y4iWKwb8ENgXnBSIoQFxTGvvkT
WFwwRrxhHgWzMlEGAl5ue+1x5rOfErEFynQ9q8K7un+9QaPDtx8271h6SrC5uxm9
mzB+2rZLOE6iytalSinYYX4CrLt+yPLSw6FqXD10Ias8cnRjCO3PpPGVsPRLfbau
T3karyPcPBLq31v1DqANvv1jICKuNpYuJlZhsGtbTDwrx1/Bwk+Bh4hd5oFdVyGl
bpz9p/ACIsq9VyVhQVNYButzEnyQxM42EJHzNBb65P/YCHPge5xIFxBa/mVEAyv+
8dENDGNIQO2siGdMzA5STDvuhFcW8xy5HkGxNBDJDNdJD7gRb1hvcxKo0St1gghF
gqkSbYRfEAnxyFCaiN7IUyrnHQy804iSufMw5w5CnTj1IsvVKBIHtS/VYfI0dUqz
3HSA8+bJxTrkJJRUnaZQskpGHUJZhwFZVdjYLteMenIdeZCegYXba7MT7rWAG0b4
SGTefDNkWozA+9cDxakCs+CPV9BDnkQLJhx1VOTiJimlw/iUFqwo63Ppz/+vwAAq
RRbWfLYjmFHXaUFj/z7jut40NGbpMj5z8J0LpwHiQ1d4HeGM1JdnDI2VDEOM2BYr
0kuFsuNFiulzOffEI0z5XeIkxbOje5L1zxnem1zPT+Y0XXNe28+c9oFCk9Uvwc4v
kEDAujw1n7hgQoL6DKaXlx+RIhRc2MXr55zp+M8lEek/2G0/rweMszIOwgyMoU5r
8hwyWVzcb/IHsiG4HHEXbW+9YP03XayoIRc/Y+vuNCgucib3E6eGfgYaNIC4QhNo
Zja6j7yCJS/egVoujU1H8QpaEhH5n5v26GiT+w+COxlBKUPvtQ3r5jBaU5z9NONi
5vcL4+60BKXZtFdPR7niRYB/npDjbgetHFv9xtvTT7SjrHwKHV4+q8xlyMc6Eqtf
v8BUbDvmewKYf0/wf1ApwJorMLPfM2O8lisVmb9qWmrRRiszEgwamcL71iyUuuiu
KNIby5VeSgtOuK5RaRFnkrgjUMKjnBcgS1ByxIJdKP76lVQsKRkntW5rTwtX7G8I
tWA1l9yCidszNmCvsxpELUbEEtjkEoGAMchbke5IHz6yq44U/LUTNAgLVvU1ko+s
PYpl8QSld1SiL1xZPjJr7cVyDUnZmG8J9c96AnLa0uNRBsja92l12wwQfD4XX25L
W5CgThHLhNPwJAFOBS1vM8SwuJJFcZWggWU08oURpv+MXGHrC8wt73H1/gpUO0em
ogin99AXgPhFFJz/iAGu6Vv7Ck5yaxhILSb3ABGcVtHvByZxqAs6Oz8FlJy1/0iz
Yp4seghI0lOziMEPIviNVjeJFHs7iQiusNpIGO4hggOilbgf0Utz9cketJa0uxdo
YiFIvnrgFvKdsJzv9DlFkUNUdf7OnWA4joikzq1uwXjN8PATaFwdBR+rFlpsBGOR
C67xhVXEnpY9ZyJz4Q/jPEQoNolVf7vlv8gydtYIoBUqwBaZECIwqDhuZq/5LKo3
QV8E3vv8j+Xc5pXxjZALz34JNtjvTg/yHodyNXPoa8F9GibAN5C0yGwa16hXBN8D
BJJrXhXZnE7d1YBw7c8T20FdtPyqgn2PLML12rT+RwB6lfehkumSV/+sOdMf+p/0
xrB2rU+NTCkoIB8Bxz+ANAZq2NmV7PfX3zFsX0IW9zEsmhZRKXLym7hq/DDhTb0R
z42jqAXoNDfG6p4uW4kqa5nQqDo4cBrjGQuOp2BasE19g0/1CVUjPf/rAGyM9y07
Ik/yWRGsje6cBYvUKA5ELm3A/WXbZCJ7TP0Bn/m49uGMA6DzeQCKsRS+fWJKIa7n
1kbxmX5MnzeV/bK4PWJoAon481hRvqA8MRhqxMIFelKJtwbhtk+dBFvbTBUG/ig8
cZV8uU05dO6CicjvMWZIHKhtG5b2rpGpaks1fRhS+H2LpODwNwQTFOeQDhnvzHDw
VC39O3UMEp7XcXoS8jwLeXqIh78bM2u2O/jNE6nybjKW9wYDOM25G5A8rxDZkfp6
RY6JIYXkn1Pz5FzuqWwe/jqGoE9v+y46vfkd1BArbUQXeIrZMw0AxsvIuJ49hkD5
TprHiXuHTte58J7ss6u5y5A0whMOo0qUCjBmNRM6w7Co/qNzS8xEgTM3bPKRYmFJ
9wtNy2imtZwJWEsMklKgZqXlzQNioOEU5B1b92wmlwF/YEBqDy1bQixyZkGRbcL2
Abt8h0gObOxLVHRNG2JOoNjdeqsOpc+ABuuVl/Lv9+Nf1vxl08KYhGxllpSMpMPG
afyWf5dnNw/PTY2AFBMqgl6YMNIsnhenYNOosSLkgHKfvkOREj7FAbADbqCpOvrS
3ZHFTLzBXcZFeDZf9cYc91OagLwLW6EZT2g6TG4ghURquEd1Qy/vAkRrQHrsyZym
VaW+uq1DHrqHDtqd3gTFst/cIScG+Pa5+rdynBb39iXXHkfpipxq4nYq0cW0CzYI
6I9wnVBOxn5ug/lUhOJWz1+cF1BZNGVBtweWggJ3kpgVZfV7NAEgf3RNF9XSDhrR
zxzw/kK0WMxsDDGzQyhMw/hp5hBbgkSG6QnFp2VYVEOczjDE0IZDnPKldi62coJd
Pve+slb+2mzQFHaQH68pjuWLRPEq7DNO9MVzwC8OSEYNzaxPQYPIMHEvvYVblAHI
V3V/qS3s+mcdbSKhXBhlGxLkCcKstUA+11e7veZpOEG1sObqnQEy9kLBFzeb+GgJ
/k9DmW6VzaUBpsT/heTL2axxJSoT9lR9l20q5sEcpQKnFfv2mSFW6+ndmZHjpuM5
WXvli6jGrKXvwd1bFdUbJHM2nAP2N5okZa562xSTBffTPu5ikEB0Vf1wnx7g1E1Q
uAa9M98JEw+0l8sWoDr7UMbJu0Hn4G62SV3TvHUcAhtlNYoPVUisjGrwsFlBZeJ9
7zKhAEwujAH91juh9ir7YKx+o/FV5OsSEcdSOa8COxa/0cvjriUd8Un3YwyWwQ8L
nUPRbX6mN83lK7yENRDZx4EBKapgVbrcxF97y9shGnl4hkNg4UEx+Q5AOmXs887p
lROtDZsyPc41y3LYKhjvvJKOxu93QIHom9nIcDsML4rOVAyfaq7FlrjvXo+1/tHi
e36WrlKvxkd7/4k7LAA7fA2ZgBNQJVA2LU5PtXBiRY+GylCHmi1x/oyDHS1ZaYIg
OniMXDXTNtMJlvYJopUunD0x7ih3InT+U0jWs8k3efMcOYm9x7UlxBa5qGgMOqT4
PMhCxhvbeVcop/5QKQBcIksf9rbAxKV8V0OnpFu2ZVUMmrADwu0LYjcFuT7cucOP
wqlYdzGlv9kYQiU0POCnN8ad/CDqiWnBXmPpGcncN7ZDFWDgll6Lh2deCGuCJcMI
D2aBL+JAMYGMy/ceiH4S2jx3Qq4c5irkzbbbNQldZ4PJct2ePdScctje0HF1khfS
b82nZ7WlxoooBDRuKPjTGHVNxFcacFWuD2T0fpy6faP8bq4H3ruJDmtjKKljF+/u
AaePBGBB18bT18gGdrfvWj1fIK0ASVrlB9NOnVAutaPWwdAqiS5GA9jxTdmR/e34
sF9D/tgoCPYwZT0uB3UDvFuXEQNhJP0hiudY27aqAk2MqLJMSr8zI/l4dpZzKiD9
mzG1ZWI6X4ihiO1u7NGZtjjNHfOUZOEyXKCA/h2JRXF6JGuYuQLEuUxkKWVJSXOB
qu8h2nfbb+UkVAjan8+cCvKK24s2SPOGhWBkJj8u2yzl9Y/8qj3UEvMFYzLsF922
0U/fgY0i/zrd7/7mkSjkZHfJKLwpc3sENG9o5ziwbGL0KSDI0Lz2sDsarciQgs3N
VUVK1dgZb3FAte2TyXMk8wKJBo2sWQ3jXss3Nla5sKlKLe0iOT5R5KMIaLO6TAEy
tS2fxDEsjYYfYtjc6VSZvrX7ZXhMNou3Hx1oUpLLCQcB1vFhOMUpeWBG7ZPwmzYk
kE9Fe4tKVFt6TpWjeEqR3Z83x7fBojFqk3VgVS7h++n478AiuvUZ41653VviKLc2
K4+95KrZxtjk14ytKWFJhCIFpUPb2PyWrYDIVFDziwGLGWbT73ESEIpePR0pCUD/
/48FuKFYpLxxKPSZOoF3DcalleMFiDnZPOVp1l4RSi+U/1R37dPWD2L7W0TdIdLW
w6UHPZY2cmuyHdAmVoeBzRn4C3j3kz+mkk3E6sZkRakvt4DrxG1c2TufqhkLQ7ee
dS0w9YS44p0AUXjmn/GEWDKjRxfrAuk970iIUeRA1KrIaXtfMSxL7MxxTLYVAGaG
JGHyDRQgovq4GUrZWYjWElPlhWFB7obsP/xYlbIV/eE6LSANK+GzDWg5aeIo1x/c
/6Ws1Y/UJ+j5gpJODdWk04LDKpEeRDDPzOq/fj4qVKHqtxB6cxY+eXa00L86dpMn
j1s3izpdn2GUJnGfFDe68ogevqga2wStRtRNIBzFhEQBQ+1s5+GZ7xU3TOoI6UTo
+1PcgvgM6Trb3wegrwhDTGldfyiFXIAXrdTe2CmeyII7XbnowBHtrlp2GkbEdzin
cPJ7mOHVMH283rMxAhvWamSzsnpw6+aZsCITeL5kJoJXmeAw1VbH5Qf/zIAI34xH
tV5ic8RBlRMdf0ZRL6dp7Z9oltyFaSIQgBUyeDM+su6VPMn7iXWuX6vIKqoA2Nw4
qU/qN4AZ9WP6++0z2i1j1CjMZDnKSB73MBAN1OUq1EBditVMdX8bj+FGfOrdSMr6
XB4M7hRhtv+2dBnvYq6ZyS5CfjkO5gY7WGHotRQfTpo+DPDYPwPyVzOOdFMmGgN8
zcMlH0k/Ynkh5tz6B+BGvkHPqbnND2XXz3SpSZgqGGyVmbZ0OcpiUKTP90itfoCt
l5Iz6D4tPtL/V+wPMLfXxGN846FNs05cz5HMWOzDn2YNjvvkgEAUVdvYNChfaLjF
Qs8L/JVIAb1Zp8s+YH45e9uvTv6pslOQ3UfaJ1wRpCrGKSd0EGgYZo1FhUqA4tAd
DLSdGUkscrxmv9G0R0BPq4gglV4VRExEYotMoEx1DAc7AJHAfp5MOD47iEeCruKr
M7NFELq4P3WneyrtEjXiGQQzsmSRhfCN6BpDfWNZEeiIj1qJX3rDTw9NPhWgUo8Y
5iA5gy5lhcgMKgw8IJP0xAOxFWUpPiQU6YlCBGp32NEvleFEntwFGtkIBJQSnxyG
LsO3pzLqH6WQW9YJrxqcB+exgpOCEHBJUM9O0KwFJeDXpxiIp3rBf2Y8X1DprmAz
hszmaDF4vMjD7Ke5yZPHgIrXREY2QXyBwnCIzDcD0qryE7QrWvoD5aIVobemAVYe
r2Nt0HmEO8kBMWTg8sdR68nPl2HsN6DuDczbhcIooUPEqzIZlzvzevNDgLL0LVZM
wALe2OY7ZG+fXGkap9Llv098cgO97jN3NThyFZ/cgM8wtAv+P1IFg5dYcLm2/uQJ
4F6dX5MHDrlO6HDIjunldTQneaEB+XwbwznNjPCyZt9Z6UDbM5L5yPrWVwjbxuxO
CeNuORsQl6pLUBixzTstd1Y+aZqewgMePOLu6nbJM9NkkIkla5xCgJXm6LNFtCny
9hyZG7+OuMgR7XtrzhMsQD4bsx0jopgeWMxz2vIECCfsxf1Ez+DV7VlfghaR4PP2
EO26paBEMITnpaSc1/Q5ociE5Ul0mXpdnE7PYWyzOo+RGt7CYEd95uEFiD1oM5zD
2mmkpxcf4PhwWmnzIIZk/WJ/tv9Bn2HJdd59LnXE2k0zWUCOX7jJ7ro4zjKZlCJd
WI0890Vp9aB4TlVwgQ/zdccZu1rJ8Hzr5PY3ZQRjX6Ve4ndB/E6dPt02a+5ZldKh
krt7Oyx3dNdu7w25DDaQTsm3Qhv9xtUi0p37DsMBYPv1pcro2dtccRgayzo+VwOJ
qVn5Op2Ztr2wWsoyD2Zoqg3jatSFr0p11NBIiA/Wx2A7lXJPUmwSDNcz/nAzYok9
VrJY07/PWnQSowNXWwn+XKEj5HVF135gqv8J2L6vrBPMzfSbrgaCr18QdVPB926L
pWH3gQmfjjM6hk3j8Ec42wrgsbWGwvvKlG1N+HUwU7It207McJeuWTYU3WvuQl4e
J+QWn8E+o2gPtVRTTaDhkWxZ938uV4KZ7ZoopNWpopASiKK3Jyxy5ziSsoR9Izkb
mtke8MuB7gHUZ9LVXiukHuot8xzVJFBUDD6/FoTFA5+SoLailHgkMBTIktydGN3A
Q62JIVp/o6ifh4udgAVxN9PeQRFedrXIqEoFajywGKuT8j1UOz/UJE1k4kzs3YA1
XxC+PGjj68x2A3tXTnyW2WJa0UXWBE5dbYCqn8zpbITJAfQoS6S5xxgP0Ezg1LUA
Q77lGHQK+EuSeoqpLV149OFK/5i92rfApfyFFlP0GA3dvdwrSPpOL0OcEsXEL46b
a4mFJaNpd53CYexuH7H0vWfzVzxSX4JPE+lgO0sq1wOplPAHWfVLUH8EQ45ioYoH
P5sWoif/MHwenp6dnuzvwNgZpqYHJZbYQnRt2HQYVcnvGKXwFm0tXzhzXYlSAFS2
GQHTA8XixP3cGUnFRABJCNDcFWWpcy2GL20Q2mj1UcB0mimSi8HEvIPp1FZooSCj
xRAgu+/DTtpNuWfHxqNUpu6Y8HvlSIuqk0T2k89iky0jYHozDyKx0sQWpr5vFEHG
SxgI4Bx1aeNhtvq1K/MayDlqiaB0W6N2CjuausVZnt8JWJM/8RjvSklqzbeMgqiR
eUGBpdgPvkPT54fAamgRKc1i/DPPomAAEsiEJAGYAsjXWVGgmONq8KscKXNkIVi6
Ur84DmxKeeQ0Joj2xPxteY4zB/5XyI3M0ctUgIcLzsToQxqsmf/gOKlF1cLC/ofQ
vJPH/CCi3pNmciKc1Io2etMcJ+MAqRgFtyXB1wdDad1fCHiiLlbwFEc9yxUUDyxI
lzBfQUBl/v+ASJA2pbtqxqTGjB3FnjpYtM28wkunUYt9mbhya8LCtXNFdPxEq4ug
j/x7UbVnQLmif4uRYV59XyLRpxipJIwq9Z0Vm4tTfHpaSwDgr4OMjYOZFlxJeiv0
qUx2C0TNLFt0Ic2QNtH/O8KiduzZFc4uju024E+3Gh6CjxVRSvlJ2OxMUf8+pj/V
m2XBV9GbeMbxkOKN7OFrG97f9wi2vhtnxpCgnDu66YImLHirQz5sQuOdrVLY3jq8
Zea0yNU+SHzIzdTAd5o+80U4B6g8Q72CA1/OgQtXc19JkFoW91Aj/MnHHvSMvOnh
itaikKRnzELgDLJc7NSrHtrchsW1/S9RFW25FjhL02rgw1eJf3Fcvgu5TGG0Jb6H
RoJglUbicETqJeCEgPHYwWPxJ4OxT0Vbo96LEeRA8FX3UHtsLsmpw3x4tqVVV/Mr
NU2R9uhy2a/aJ8jKscQdu3pIwBxsPMRcQ35skEC9ZGqH1AacvM9vylUyIg5NRL+b
sRfVLtKhwBGG8FfujPJfFGhvi+zSCWb/bySeB88wRtY6wljUok70VRLEYnTDFTTI
3/l7VKTBUauhEMWC5yw6o1ta7HBzn7srOmGTEmbJt41BtOmmg+eL4Y0HwnAmv4RN
nn40/z/a08rz+QJkWnuMwbyH8g6Tw5ReB4YeNrPv03nO1eY82g0sFteIAir+Mx7Z
5CbK5vtEtkpVianl7PE9d8g2YdX3rchusggT5xs3+/R1DLrKyF0iQHLLGfZheub3
9LPEmtpAS8uXvmSuioy9wMxpjlK9z8ez1DueduPcFFl1E2YCRBX8zNJn+W4hiamx
+Tos3wLetwq790rWX2GyuRPQRCaC3S0Xp+2OfADMgy6NsVTQcvdLu3ndXvJd4CTy
IWjPbhfY5lgmpqVk3B6XdFVJEZkuxvSVqph5vzTSHcGRFe4hguh+QH81xL4b/yit
7wslxBJKNbXNAypqWROeAm4S2hyR8+1KVgjPWbo969oiaqD+9cm6qA6MzqXu1dQ7
HiCHevPUomhVqsIlMWhsKux5iy4HjP/nP0h6Tt3+WfvzqnSsPmAQZAayy7gg0Z/a
36VEfZtM4/sasBcQDvkii7sLAoUcuCisAUr5uB5mAnpEPXdzbZ465dvSqBy8XuLV
WO/hYWh9c1Cjs1qkuXoqbPNiVMofMM1Gg2fhtlbZRt6o7NGPOZjQ8785M1fOowcX
jzT76kH/wH92GauFIZ/Q9y6hgTjq2fLTEYz1KtJyzzZg9VVtrOzAzdhh/3/aVFvS
wvc9F1CbLoqbwzEbWyPKn67Ie7XWNy0pT0LE/cfVaXrn0N1j9hHMfvbup6M3ebPO
Y1uLi5ddoDf1181UK5tS8xdTnvak/CLr3eee41oHeYrFFWzaaEwq9C1sAzlWtgWJ
pHTyUcC6ZGNS4jX4qHnirWS1/QjPCW2E1KnYBdGaclJZhg+2jKpmmZIi1sy5hKtK
A5OqdVcjinFKS4G9SLWkwhEC5REeFZEqXdsVHvQ6zGiMhr9pIwNXILhpsI2Zg61U
MtpAtDkX7lPutCvwWINSSNn3mVjyJSDFmRQQn3sPZxS8+4ghi5aYjgNuLYXRmRvg
NQCUWSQmVj1jmmRIwLlYBlpaO+CqFxmTltIcL6iW3OEp0SUu5UXid5+oGdT5mzs+
79z1Eh2fGQEDIylaIOPX4lFc4ZmoH3kFc4aUX5IIf2hS9jS9V4umm0uk/9RdnR+1
HF4lUHnBYt1YIb+Nv0dU4SC8XQ2diAst4CPKcfmApKmJTSnu1gx2DCqrvUtwwCIp
G+fv/qTaqnI8Z3SS3DHyE2F1IN7MfcgdNuGUnVc2NIDFeyH+9RH7PtvLJmAKJlWc
V9kBA2o2W61yOGUGMFkOgNjasBFhkkvAVtIi/P35vdzChhPRICzDnEYkxYcX9mgN
tlWGpDQQbBS55pLjRYRJbDazIAPfLs1DwPELVosm3xmZ+jOik8clHaiyw631USyR
jkqukpwk1vaZ6IK69ZZ6tHUy5Yid6lApNYgj95zey6cx1TVNq83iXfUlCgniMmqu
kqkZvcPrLQVJszLXGRJe1ueo74BEgYEpcGBANyubJfJ05PmuvMPiKDUCgKsTVusI
4dX0PtE/QqlwXvMRCkCCFzc8FW/yzDhlDYqz4NVPM+GuU0b2CU/yUAxAz9+ZQtoQ
aktmjJBFhVk88haBAI6RwbQaY7k7VN2nInO7XNfVw9ZarBlS5TWeEOFaD3zUuvjw
CLLvIJYaLZrPTrh0KIPyi6BiRBBXeMewGlFm9pSuRwyTUbqq/dk1fzasHZe9Vthk
/L+FvMo5Tfqi0to35jnKFi7RKHH/9vM57tXE/I7MuK4x1WiYMjT0VLd89lBFsaLC
T52zJm6YeAtLcmcqVivUtIaL8mL7CWhMBg6wqC4m0L5rpO+6yfKhtXvnzk3RGOu0
fKbDDNplceBDrVG0QzyfM/nfscoy/M0XzfL/OOHch+sro+K0Drgep3WNWzlY/aYF
Q4ugupGYywEYZayXHJ2Y0IlJx0jFy3qG9GwpfMJlWbN2lGJRcboEgSUeu38n75dW
7JCxM0nsHTj6PhQn6HaeYqmb0s/vpbQ996OX8EkdfRM5hFm13y2a1K+/8FtTUrMs
6ZtF6khU4BHwqKBIh5FjO+4/RsCUGt0ABqJa8cCOflhx3zJyMlTtz+XWRxutGytg
SReYiwMmmjgOX6KRcfAr5mWSdXww35n0WPcjTq+jV9ooYI19tYhqd2kzdbSIimC+
EulnvBvOBcit/zDu435T71t2eBuOB068WWW5wRzJhPB+mPNouKCOJqY4+Jki2Sa3
HMeg5oSf2xIDEqAXiilLPJBCdPfIoNthZLL3WHhF69Bcy8VbTPklvWGL4V2jG8+j
FVsIJ007lHnoXlYzd8DCTM8rRmdOiPNoBhIk83I/b9lK9JkR+RNvWPEm/I/P8tTe
EzyYIIqY9Gkd7q17l+yebFWeahXCLyq9JI9yPTcohe7dnbpNoDqpdGgQIXK9Q3pQ
BTHATDnupwI6FvkUUJXElE3vf/8KpOUhPLbACmmP3H3ZUKldTTawfEgv+SvLotbF
VM0BYoWhAi5MZwR7LCpej3l5pDWVwwTuOe35A35VZYZmllc2rnMwzO2SV/fF5dRs
v9RiEsb5G49gObIq6urxSbR8Mr3sqFY/m+PWW1HZO8pQw11WuQqOsXK1rdmROp3B
dAxA1xvEQ5c0jdIRS0Fgmu7MmoLoR6qoshk3nN8yPwMBubqh8h15UZTo5wUAgvvY
2q5Y3FaaXK1UB6fwdYSiFAJNeGwtyXgiTscDamqjrUyy9I1p7SrY/H5IYq9iOw1s
j6xMRGBksFUgnxGj7vAigQAjRAKmFG/ue9Tp0czG231U+z3pZvXZQ7Vm0jMDltU0
g2QzWlSj1opQLseSZVj1Vd5nU7MSnr4EsbNDuvx+w3XPhB3xEtIgfZb4L3K7nSrf
MDgtOaXh0ATIspa1rm1tYGJs6OlGCjLWPGh02fRsQTNrYgcuBpAAe3PFUM7uvyPl
rxkMOjNyyZ0paH4HRkENjfB3LbxrV8JI69/NOj8Aocu0fRjSBKrZ4WUvs0vH2omk
odIK2FtmdiqpHyE3Be/HD0VhTxxsk7Lga/ec/DHJ/7+g1Myg4Vcfp57hUQTN+4RA
yfFELwDdkCAnaFXqoCIwslUObbtjt9NEFHsb02fRAtPaySRkzz3ik9Wzr1f9O5A1
2hWs+LF9cFXMziVjo+DLUm2pyURrNOzfGx70G42PPwckhuL/NsCno6ddT/qtI5hL
kp3B3kYSqq4Blyb3Zo4hZCxJcHGkw1mCehKKPOKaVE0rc8nGg7SlHLXcl5VxBc/W
AF0mQwTN9S3PXXxFalTYnNc+TJfB/IGybUc0F0a/BUP01xIwCBRoGCmRR06zTiB6
abM8f06eBi8b51BAo4tn1pY7+LPedaeIsR+/Kl0sqUBae4EnWSL25utRIyooIGWQ
N7bi/GkffDsl6/w00tQhnxz4kWxUX5Xr0LHkqD0SgvjriPdd1YFKpsM7ia1Pik37
CGNvauWlzATzd1mGhXIn/RRtZY9MJ6px2hso8++ZgkV9mdhJvlKqLO34Naa88YqY
+QwMndG3cvcFlDGE6yIY/OwKKux6aTKSlPNLOpB367grq3lCdXop15qct13bui52
yScljByS/w6KGJ9q4NnLMbYAgtFNCuKuFwrP979eMLSrHeq6emGcJi528sAz9WWt
CH93PyRCw8+/U3UxD/quEFTFsBFvGpa/qmeQCeSm/Y1BSy2cUUNj5H4/TUA4vaHJ
ZftnlvYpQ+EuhvkXkwLEBminV69cpPBetEpqLZ/+e22hV7lkVYi/8AQCijannMuj
pjjvqqdBEB0uRqlJJEwUahnMkihVBian2B00/W6rriqEez3nrezsWqwj0UHDoGeW
XGIrSZL2oghzqGwv+jCs1xEPqddkIi+IvK75rTQ0/gQIpWMRt8iNvxw+RQmLFoL0
nTOPWs4/17koNgqYqWxBm+AzZ7VMRgS+1Wfj7f65mUV6Kf5T6FN+MZeWuhI4TXX2
I3JmqDsDP9C7tYFh+LTTKU6Leg+kBVdFn2T/tA8HvDPWZG5I1JDu6iuSV2ogjee6
3DhEwZzEcaouuzxiIAqoiAcABzoax+n774hxVd+llZI1PNsx2UvAOOCKDyQi7OOu
qZ+mpqgHWqC5Mujqcjm2Qyhd37z/nD9AcmQRukwVIC7INQEU86v3NxuHoOfNXET7
+nNRWLsRzDhdBqQrWmH1XNiPUXNBRb0v8K6AO/cJy8DpUbIUcYhM8yZ7MpkWYLII
m+O2FrtCk7Cqe4wRo6opSW2MhD20FjsTc5lNLMJ+4Rwiq+7gGcEGfd0Gn6/wvDCt
vZmmfmx+1GjuYDIXQWnww5uH7h8dis2Bq1DR8c4FS7llM9i161DWXCPaW2ktCuVh
6TsXRFgMh6NXpWHcFMThHHbiFh5e6fbfm25nOjdAZPktx2v0l0MyqcuSRQyZBFY1
sva3B+FH5zcAGwvu2V99xCyuQD/H3/WDn4rlY5odZhAK9bOG6akyRlu1UUExLuOW
1Pa91joA3OQh9uISEZG3Wm5btn2nmQp1UdHZzzZLP7SyJ+aPdE4RtmsQenyY6rtP
dS7fhEONAiUAeIiM9GXs5VpLv1TbqaubPtA7kXDv1E1MBfT9K5m0HbDoRqJ4+5a6
ADQ9HiW8OxBQ1fZlt0UKwmJgli5FcmDooYdMG7TpScvhvAfbTUWBQfh9wPo0/Uhm
JG1W2M4ahBzg9RlboVDwBOvBSyXtJOMZWXQW6alsQnilUNOmcW/cbDkAF9Cu49+p
8GQKkthYqXrCQJjYLe7u7CjJhisXFlLRC6KDuy9pkjvII9t5Xr6SV5hFolQDk4ja
5ax0d2dA1is6mIKwq2bg9uNRgC1s8b0J58xj8TwVUCyZmgxQ1nvkjxMLefGQn8+y
MhLZXXyFWCJ2OkZAeU10zZikeX1VedpdQPZuPAVWw0HZWmz+jc6i+2jqZ/rd1WIZ
FB3ToMTacTE4ykZcVIwdpZk3Bo+ygidtZC48przQhetXk45PdZxDlDmeafIlv4K/
QPnfEaZVG59Nc7KWtW1IRcL8HqjaWKL6Tn5QfevJV2ghfH/43LWq4APSM7LQqAvV
rwBdMikH5WbqNy/D7QR3A1pz4rFX72x/9UPT0XJF/3gB0hM1qxlStm2kKcHxZdBS
CBYhRSGeEoGoT/Khz/O9V6Q2JiKYbOZGX9jbveiNvCrZjTBIvd2ramZOR9vjDCR7
uprUybwP66SJCxn/YRgFr3W8LP7v2amheFgrUa5ixnegGyCRIX+416AMNiDicSeV
7fHTHTmX4k58kH70GSzMUQIYfqKCIy80VC3FN+cSxRbxUWzTKY0ycfyQ7VSGPSXf
mRGyNIgjkHsMsiw9VKLp/ndOtTj+jKCtN7Rp6/QEUCcjU1qKuiimW501b7quKhLN
iSEoz+U8aXPF62VC8BK5Qd+W43w/yrj+/C5IiKSF9TZPM/GhPzrEvhlJy3W6ClNZ
Z2m8NosmLDM1CbamAylRmYuhZORezX8rFbeWNag32FUbEVCc5cJZRqrz82jYn22p
00MTYaSgfXvxXOuw/VA/DUXf+hsCnp2iTOL82/sDkjUqZPC0nTGNfxj2ZOIDwfo4
5cYHczGp3BtweceXdTAY92unUhcB7OVK84ZT1hXmTNzAw0qIkAtOyWg79eRtSV1/
dG/6aW5kUz5luNzkBf/dXwSrFJW0zTdu544ShAlzjF7uhQ18+Wwv64g21B/RjWTy
16PYsjjqzlJ6upI68MoANUtRal3V5AvsTt3OnQQvBVeUI/F35ZE7UfpbbbPxCLsp
Pev+TjcaQtvCOZNblUTvyNMjSI+n9SQyABZTse/dp6lmkzGl+oyyQ4g9yPeRHWK7
DXsp2BsinNS6wd5/ph0CNsLr+Qg+7B9ZW/CKQi+q8T317fcLd9o8t48gj9jxAc4g
aNtonLLxDC2EZP2S4ZfT+3QcqaMpGxCgK58TNTFj4wi3y3YwjFSFVbrgnjmPwZsP
Tu0iKVAMXnuudBuoyr8lT8wndC8bpV+SA3CB0wkxptHFXSEa9Y9pyNCR1YRPpRGE
Snv6yMQ2QUCNtkQVOHHfoYbXiRHUdCOnC8xswseErUe1Cmm1sk9ERw/bO4kTzcKK
D6DWrQ5BpEnnKNcMAryOAlV5RMdayG6ksbuHADwYhMuzbzS7zAYbvGvMQgcWvitv
2RC+nRK9wD/y108lCtdJCcvg6pdMSkTnSfRfuGH0A9aR85cgCMehPIWy3gDD2k4d
MytU2kU+G0MN0VI6FdZLzPHtzpWDWJa3r1cJE6FmdOYQ97vpuKf7KBCBwPx4AqMo
nkwwyZSPlmKyxWCaE5yD2wQJqHmxfy/tHfj1j4XXQIXnwIgc6CBc/Qwt4NM/BZK2
DgzPdJXCk4p0ZDC27Oh9pgUry+83SV8hixQkDsHWQRDJQOG4K9HhTN1lP+nVX5Vo
ons+ivwIuUXrRnCNcWjnqYUs8bEVclrf4/oqWOPnYOIOMKCRmuQIiZVfdS+gTr+S
nQmTvlYOqIDpJoEhUKa7NlRAjHGsQvPx3vT/a+VjxLFnodA+pE0gYpFr2mNbdVZp
VYcz8sXFe6jLLoxV6GsNbnPebcYgWH3Z1VN84d8De50rUFTm2S+Yl/yLf8wZDRa4
FjCRRfqDWGEmzD7p0FWdMtRp/morb2eJHDtmepLihj3yQVVYDZ5+pfF+sXOkFfaS
jAfXxZKN8zTc526dwuxfx6JWYtPQaXGc2RB8jmw2pb6VS61t6Ay0Bebp+deZ/Tpl
SkW3Om9/6AX0B/2/GpGd1HxFFX9zu3S3QUX3neJ0Ii7GqTDtTs0cpWHPNk9BrBJB
i9dytIaPruarxdzRB4DqTtVRw1p1lQcNGybaUgOlqa8bNfC4NP6WODPoYWQNqBB8
o8ubNs6Z6DOMWCziOh9gFt7qhEWCATylzG1IRz6rAJFewGDe/3Mvsim3wHWjhIOO
FVpvOLOOZIYJ/8q55hvpUd9ZOLLMsajDrwn5hQP1f9dqL93u/i81Lr4hmoGoYyoh
ikzHqZiKUpBt9xGUBR3x70iKZ0awlPfitbsiKLwenNLQ9zzF59jOuRV5RaU5SYuu
dElm/Q05widZaGgULazm3g16NfCAmVRTj69fBcBQNx+MNsoZJFVKcbE7TTgm8TJY
C8D6SE2+fKr3N9ldNWj+1dCYF5JxF0+LRLosGbwdZouj7YU8StUKsm9ovnGhzkla
e5tZpVbAwrZhxQK24UA9SazFGPxIjxVuWl5Fi9bRDTOIMleQ3V5sre4fYBE6XcaL
itmJicu6QX6x3wmtRar3IZ/iDcGHZ09uj98uCY55it0KZCKFaR1LkGGCympOJ4pH
jG5krYmBOZifPUGdSXSJXYd15V4H7UJSNXCUw+3t8whnLQrhV2FszSafTm94v7fS
D+AJ1wiqdb+IyIEb6Tk5nFiM/OA3H2Zq6S4km3df0fbVKdOHa2w72nrOx4nyqfjB
TXYgOVwE1AkEmiPGmM5wRxoiFAAfQutYwkAW2PB4plI3cbUisv97FKpSUncmG2oR
5uSYGq0mhzG3NoV2AZMaVLII6TV37h/8ovQlUqrBERYBhZDVS+nrW4cRXIbfz0b6
1kS7zHGvKKW2um2jdXATYIbxE9VctBQswpg+b2z/j0l5LsTJvMxcH5MuMMl5143p
3flurMQ5wivkGMR5GLkXltuML/xhGI+RYqt7UhQvVF8RHOOGtOoh7pesGrNVhZsW
IEoOmK2DNSQ5PICHTMXRwmjUNgCXbE1NcvQkVbvnsbjaeLtxfr16fqQOIic8RMfR
XhJx7+NQTxCwLXH5/qUV1v/Tf43jbOPXrh1iSrGZUk+5gwVb3FY2TgDBhN63aBK7
hBTmzwDAnJ/6x/03r4YF8fQyXlC2FuD0S8Wyt5bzxEYTa8m9HQ+Jp8rxeP01N65f
YqZL2pcCJph4a5fzYnTMAK+lvjQ9pqXlgM5KpTJY+Et8kckTJL5gD4DyF3vYAPgD
mOmoUPeg8jOWZQtFTOcDo4ei+Eq1+R9q3mJ2CXrmxbwNsMbYPN/2LBLe3EVkIDO8
xrQ604z/d6NC3M1cjXopFiMGP7kRyMD+Sk7pE+3En7dAdBuhxFckSaTHaSfoBmX9
i/ZYM+QaBTQHzAIxBpjlRGf0UZDC0l/dKD06He6MIJqnlhQymObZW9YPby05DU5X
0+q5g/EH65+YfAMwuX1Yr45MXvgxoMNmYN66zDKGD94B+d5D/B8+Aq+7ydesJGZX
k8Poobc4LfBND1c8pUNbq3sryR6qFAMSioDJB18wMJ0Ii5+8czmzP8gMvFyYO4SK
tMTTIxyxfI+jZMhnofvzMhY2z8/3l24PxwswvRRJar6BGLf/5RwVu7SVAi4M77ao
hNieqmfN81YAIpidhJKBQkE9TGt4l15jqc+g7BKiKLhRyb/AQ46UJNmwHGMMj7lC
Y2hJyKOEhCxjpwm8MZeur1AS3wyq1ZYXQJrB2NowNpSSbbBKLCNgt5vEMrHyjwNo
uWLlADSoIvE1/6UFoxteR2QZeMh/Oq/179xJOOuGHDx1EBbwrYSk1tmRxKvITw0D
BmqcChfMSbi6pK09slS/p8rxrWkp2YVdJoZS0Dx1CNDStMhoRWGsQpcTtwtgMHRl
feB54sShxt837U6HiwS7Pazzh9jf1K8noHlqVxOIapR7XVciktBk97hC3XD4Ff4S
W/Rb5XYCSev/2H1mJOuTZ22tkahxqGEXYEkOmkLwou16vAEHPXGKaLObXNrOnjJZ
v+yn/KdFnV/utfHabZv+hgXzyG9beXRI5WfZOmf49P4ggqZugUc+uKT+/IfgAEoG
MVYC4kbB4RVqXBsuwLs1fgq/l0Y/NrVAV1dJMV9NnVuVqVcBti1VQGpunTcrkkPp
arnKZpa9tX8aHM3NLYTSCq6/njKUhPTWozMODDeIoWUITcdqh6Qpyl30XEHlLcOn
ARk7iUfoFHzyDJ8MOosRzEMcumiCoYTY42u0PfzKNSNmLxzUvrHWAhwUepMWV5xW
QhvVuMcL8VcjuJODL7EtR+4M2VNF4OlS/Y3QIrM5pdKuM43122nmnWF9UMUtQciV
HrkwngS2QAo4gs9iVMI3YC7jPqtEl6Ov45EWVqEWxGqur5A1lWHRclGigey56DGt
J+ZWVd3MeLpzSc6jx+DFuALEIEYY54DurBn+oPo4WPSjDd4wzKyFrCGw4cmltIvB
aI/qV97PWWk1HK9PSVKq4+6Y8hMNiL1dvc3ozUhtSOlhbi6RB8Q2jeeGFC4UA010
iAczMsLVjXyb/TpliI3PLXz2uJSDvkZPNsTWmfYdjGyQf5jvK+AsQojR6g0oxkAZ
5Ok9nZmv2Egz5kDrzvs9nTwbRfvXM2W1Xrvd067wC0y2kC4t07ICatOFJ7x4i/MQ
YZxxuyhl6yHViq33SKJnR7ubTIY8SIFvsnvfCAeKwaEM6Z30uJ2qZNEo80xNnPrV
wcZBgabuhogHE5vKJj3b1dTR5bfktCB9Wn9Zb9czOeH/CnwQ+6FMGCuVvRDAGEWI
OQ8CY5Gd7ABzhst+Xmnelj6v+l8C83/HPrc8SBVGZkTSNPCj1XoI/LjAsHi6Xesl
o7tqTPA2P0xgcemftiX79GPviAgqfSetCRHg7uApBOnzaWGp1hxDWYWhmLYseXBP
wPoep6/pJ4o6Eb00Akedlg9L1Xc+oVs20/3Wdl+4KM/sLEhy+pInWgR4qIIkI9JT
2oM0FarphiFE/ZE87KFteow5DSVNRsrCXsFWUiGaI2ufNzabe7SAYgMpTFGLrR6A
UsxzK5Nk4PtDN09XKnrBPHY+1NUlNzsIJqAJJDFEEWRw3Em3mBPzOyJVbbC3r2oT
Pz/8IeFjgexst6Ziaqf770h4LyKlhyCa1lYovsnWYXnzw75Qj9BfBInMgVSIzi5p
ZcLSZIrcILwP6wVG/8QxSAj1YfVRnIfV1LqQ7hhRRc3rjcSCAfmAGX0wkMPEbdtu
i2M87AdkJHcZUF2aOCgyjRXtCH/QiJMubane1GoZF8k=
`pragma protect end_protected
