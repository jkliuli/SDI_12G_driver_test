module sys_sdi (
		input  wire  reset_reset  // reset.reset
	);
endmodule

