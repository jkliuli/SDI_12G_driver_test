`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
tYMuod4fsW1Ah85xNoWLrFrnqA7XFE2RwImt/FuDZOiNpsVw2O0DXIgY5nL6RfOh
yML7bwKMtDkCxwArbOz0ZVD00G6Tekmv3Y/zMsFQJfwpGoKYathycy0Eqk4irkfW
LMnfGvTTphLcH+vDHCV5f8xgPtsxRVzvUr51M7+o8hY=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 2992), data_block
DhJoUzPAw9XczcaotmEUWKVJ3qi1feaYwInip0x/rZT64f+6w3xzb5+kSODAjpPm
7G2JYSwKsKQ4LNSMBFqb7HuudV5OLY/MwBf/TAgRWwwXa3zDoG5BSZbo2SzIIR4D
LLzWvKXMB6Dj1lGizJEqHAHvxCoQwcMbtIF4n4g0M/d5uvF30dP56aGKqTfX1Gdv
YM3Nf9uHdf6/Inn9l93oiCHeooCxOgoV2coyUYSbJx/nYDZwQ1kjJzrSXbvrXDGI
+coiCir1E4jEkGXPxT02fheadvyCfWI++qGVx2YayfrOQSy3hgKZf+nbri4x7oO8
pAiwAxPM2Wdad5Wk24NJn10zgwubW+rMTeH3EkITVe9dkVx7AU/wSltc4bLX8+Qn
g/lu4RmOyYjlbJBBFZIBOK8RQJOzCNNFPZwVzjuvgLxM8yhch4LIbt4lvZfUEiD6
EyVPWcw2kfRsIPAvOENQoe8ME1eld3gRwUmDC/tQazDgdgMJn9p7lJzWP0ro7FPb
L/YW/UUWRSUHoI96THAldNjYMz+HufO7+rb0h57NufYBwmwlOnHxlx4+lWsW179R
dOmhNU4XXf1mLq/wREAQDUsOO33H9sGiAaUnD2qq37KwsaKKq0VvrR6JaE88/D8H
s94yy2AfIXsOZF/CoQUfdKkAJpGcdns7DZM2pKaZeb2r7A/fBRHDuxPVg98Z55lJ
zCKCO1SMbHGuHG3kg0z36BOxr4JuDV13hKu6R+D/BH4UeBRdvrBXjDEY9tZYm+bA
UacvDkoTpw6bsuEdr3aAzx+PK7R9bphPNR3RgFwcIYL9U9AJ0Nb42nmF2PKd2Bgp
5AdjbUrcAB9eSoCsxxyJeY5BaJ7D35mBJ0i3E3MYXXL5L8KBjFBV1rCdcTOC2a/A
XV7rlqKliKgWwwmA/8vavBfFKKA1tJLaBE+Jh7rI1YMwCTFV611yTm1piIinZvhq
eXDXJLSfIX7AcVlSd9lsRIYZqhJ5343TVDjMJqDE9phPyUA5uPxvcgMWXJOdv+r2
gTAWNhXucDnqSo9Zst06PNnoqIYpEYcAVBGVzXrJYObqXpNsJaFuE2nS/9w/TeKT
ITAEwUpuwLe2wv3M/kv9YLbSUqT+ASyUbRRSZK9AV4GsbqOUMafYeuSl0RyO0m8a
x+pD/vvGQpyB16bQ5XBao1dpKUXbKp2eNwoLkp4hIJkNj/32VWEwqPhevrpHOuaA
1Vccj422rv9p3uaHies9hl4agnL8zHDONBpU5uiKpY9yvvpnsUNYyhEQNgJ9DEs2
DodNQHHF4jNLBtALkapffLRtauolwSNg8kuXNomjcFTyaL0cXPptiSg9cZKi5l1o
u3eYEOYl2/+I/+6UP6JmKs2LDIjz9Mx1BPU2xlFX18sy8D3/g9mDa6Iqhf4hUNlm
6C1srdcPuIOB7K33ug1kLEqdyjnzOk0uZR9+MKu2pWGJN9Xnl+s6OFJT1uywSWk6
YyW1YhCXjB0mc9DMPFfy0zlKrbbATXRFl/hH0aAG5UJ0DOz3IXplNchIHt/gsKXD
H8S7wa0KlYTvT6tPBBcaRyX59C0z5XviOE7jtSebSQuUAtkOOES975ixJq1YjRy5
czvpjInDWrntPJab5BMYTndgaM4MO95iFR7KhlEjLyvI5w1X5DHkX3xZxF3E101K
w9o821BS3YVUXrq+Kgjtkvv3ps/4r+iKBHsIqOwTKhP3DyL7ZwXWBEUR70ymtLVU
/jUPT3je8EbmrwxFmJiSdkl7djv3ZQEj6lzKU9BQI60j2Vd+OX+1z4lN739rapw/
8hdlFZqv+To8BGaKUUHSWODltR62n7OSLI0xP0KjYVHt4jfEEk4caDnprDw3xVlI
q5Zs4ewH3h3MrTWf2qL+LMhxMZhoeGS2f/ZcMI9uZtYJQgWlNIfrj8nMPRu7yrzJ
vlhm+RhOgsEuY/jHkaeKOV8sIK6p85i2VcE0IyyUR4Onyl+am4VY+lc+o9QnCr7H
SHX82L7Sl2Ei5pbNpAtgNOoOLPqhXJHUgACItazzcikn2PptCKw+Z9Vd8HKpnhWT
w+WOM6or5azfF/8Ynklhy81QyFomyJF+/Kr0oiE++8cttAKPnYpUi5Ar6UyV1Fue
eHqiCrOrgbxo9LQVYkMSJ/eanxI4KdzisHPXBv9A50+D/OGs1XAjWRIpTMrCaHeT
Ttq3phQVV51AFYumliEfYRLg51fgIxQhyEru7vol/AeJDyLORWpVzJgcVERGvHWV
wvD5WctO92TupmaODwkHZh8ViwL3JbWuHoo05+YJTf06to9cc6N84SbNtt1izXYx
YuXtADdRx3mA0vTjNAfz2jyPIqKUd4mHuKslH+6ax/XqwL2v2jM46foral9B23CB
Ga1DRHnmUhwvzJUXUMQxx1vaYEk3zyd9MeXR0gzW0cn/MSgDyFUp8RHQZVEpgOvo
8O/bBqDcl/fRsFcpaLrmdBJzY4lDrrSIuXvIbxZ2pVQdo8gmTrMoNLeksWpuZzqC
/TCKGSEG8i5LQ05brY8mmPcd+WUal26GkJDFaL2gPva0+HmLWNTcjpPp8MGxfLxG
OP0pBlxY1Qm7FevY64+S3Zei3DN84Okp68/8aPRYW3rHMj/VRoaU/6grTHN4JqQq
U/wQzEnujVJC6XenQuGPlGS4Q27gI5qc6teCx4P0N+UtuaX8hGxuIVOvsLB43lOA
iQsbhn/JUAcW0PRrRR51ovnEFfe1B+mX13n1/fDgyV6kjdOLt2xH5mq9E37lstkh
Jd4YeQQk/LXnu8BbCTDvwofYd6DqF8sP4kBtndaG3V+BvY2edgau1byfx1t+Bri7
ohTAX+LfAXSY5eAEpVBizl06dDZ03eLx2OeZaksavs1egS7JsrnPLs7BKbfkG0cQ
wbQDKBVuuzbhD5f+dWE++LE/P8p//JB4VzW0cPcq5NdfDoz4413ReA3HMWL4TIF7
6VLt4E042V59iJPQdzrMEgllOAYTkGGCvxT85ewmTtieej61kzX7oy7MUleWy5Qe
8qz7ovi4N3jX98L2Pocwbg+b2gTRjMilZ4sAEYf+CJhzTRcyz8FXYxrHb66cceGx
vi27vCbVQUfcpbS/c72BEl7+lJ0vAdyjRk0GydK7EcNwACWa9T9e6xyY2lVX/sMo
zTsgANSoDltPwqc7mudimo+DAdN4Lm0Tr6dcC4ryUs8tKiGe8iSpzAggM7hnJZnD
CwaqhdO7fjnYBNnNXxPkn9i8QMvoXDqz6Pl43DPClEI0JZkRTWPRpQxoYZ452RK7
HQAMKNeMz0wGwHCO4UdQXQ33G5VvqC26/YW1BCs2B7HxWlLnSiN/Th33jkxGUDp6
hmQKlfm+xUf7HSkN69pWSwoEVVZDi/ozDeZ4VrZL2f43zxnF8p8giopSb51W8yuz
Gzo9lxt8rlw2MUsRRcEKiEFMkp9Sq97kt3wHE7UQozsi6fwI1McjpPy0yT78qX6K
S7jgLJNA06dmtLI38YtExpIUDRYnDyZKcTHg6AVa91M4yil0Cs1g6RTmEs/tWRmO
ErLFK4WUC+HsLtjeYYJpwiHw9EDzmOtj+I3ZFg8gGtHzNX2rUzNHqYHy3SRJpmv1
1j0fPOxqG2bMdfjG6+UJiAFCS9mVHAGtq/Xrd9Gkpj4t7bCR+vw45Xkos1dKR1Xy
JbY2h9iQVTw8F1ual/03LioNvhhY2DYrpKIuIm7HYBrg8OAcZgEvR2WLRHm2+a1Q
BWlhGWn9/IIhlt9QlTu1QK/oozxNXkBaZJaEvkh08jD9HfEZqYOwF37DhPkpkb8x
2OhM5NNjxhxoMXGiF0+i3ivLMmvBE0nui9SL+piaDMWWCQrTmy/hDPN2lZ1dh5PU
dpwPcz4DCwr8o6aEUizbQGTLBzuKeOY/SfPPBXMtxwlPAyWMI7kXs421dRFhv8rO
WomhZi1VgdeQk5ODIfi9YSRxTjTDrbHJIOgEC8VRtE056+3V9I12OMpqb2DTw1PH
zzaI6IN6SlMgO2H4G/jFnA==
`pragma protect end_protected
