`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
BbIchA/HudU4aeATvHKU5Cugkw79o7BGp1OJD2hBg6MjHUjBFauvYg4ijjqaPocm
DiBy0/7dQ4jlTAW8iTfm4pNm1SIHsioxtUqGjWlRugUXVHw9ryBi4QMgs4O3mhJh
+DJBcfQl5FiDAcp1/p0RfbJOIKXsJwO51V/yLxwq7eY=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 10528), data_block
AY3rkD0EnfR3/8OIEwiS6LGotmV33XalvZHUZe9vEQomTo++Zb1xr7b97VTcrx3v
oEOVcWpIiewkoaxbJh9lWKAVc/Hnp7Z6S85Qeq3/KrP1Nhy7XucR2CceBKx4VFLZ
1vW1wHf9P0JYhC0l99brf/cBmCYUIh8ufcSEILpaxbk5cReKugrqQ3b2VNR9A9Qb
HV/0jYJpXi5z3Amxsm/dHynIi5Y9W0PDL/NYsBJ8l8yCQuLppt95EzKCR4BYw8BD
+icCCZtIWVOHT6HzBAYANm96uXB5XQm+eyc/uUd5fTTuFEZ49+9n7hZqGSuzQ93N
1kBw8BQmIywkGtTvf9e5jI8Qtd2bENip4eosUgEbOIahGxO1nVeX7BNJBE+Kmp+y
n6ByoBQL5INK6RT+uCmFbP7Hq0D34PVBFlXTGqS5u9ivc4t5tWpfEWzmsnimP78t
ALxcuIeZl7UdHPwPt+W7PJSIxRBM6oBaNLK/ZcBoiFd6Lj8T9mNRQ/fz9Ja66IpB
H0fXMlCpcnP3+XJUYgzmKx1G8303u2+asjByVEL++UMWTfXOnC1n3gvmsuY9f7Ba
CWyWcYH4A2q0vlRzM6aEa60VSoOZRstNoXffeeLGb4DqYpAHJWqmzlP/L4BMZMdd
ythZ+IChYWHlYmvmuoOzam5Qh+sYqGp9zC+p69fi3v3DSVeOVFCudUem33+i+E0o
nG2GIE9inwoW3RMX/vX3LzZCvra3bgY/xYPX6rQ8G9mRlSaJPHpmUvJxduQ4Za2i
izO8ksS+902r6mWPBzeP5FTHCxw/jtUVRbnoUGyUewzCCBaXLRnZdqUQ0jBbVvIZ
VKFd8aJqd3ZRxr6xi+a2GJlm5XfGttTAsOPZSs20akHQ6gRTgpqlJqhSKbUMunvW
U7h4ZB1WVwyNWqrDauL/DS99Dau51fzKbrOif/BhYwAr5XZX9mc5Jlez6KM4a6+g
NGAMc6fO7+KD/sXIJ2iKhYE49zKbRspnMU31A0RD6It/pi6XfUTpQjRxyKB4l9FJ
CXKOWWw/modp0h+h/5DELB0zFMbVwIZNn1D9SxhUe5PF2Xs4LBfppFsGelXySxHl
chlN1FL50b94jROjwhQb5mpBHq8AUh5LD3WzGAQel2hg7nOuZOdErO6XVbkxNLtD
IcKE0eXLvyIhhy1kIc7ejVNyQEruQd4ea5FtOQrfw01Kg6HJjsF8QUpQUHYBzTnm
vSOeRkMhNnuTNptih1VFP+gpY/pjZrMZ4UTkcxJ6zyZ8zZIqj4t1D1aOgAvI6Ae0
FppoEiDW9nKFeR6goDyq/RyIgnYzPbMyLY/h8hZAW5O0o9JK+h0GLeW8asvTJXrR
5LjmiNiqylU7S5QfNoRCJzggAHraGHnsm9WA2RDcyAWy0TOO3S+xar+A+vazXmWr
sttK3Wkv5rUVsqLNVHGvguJWKyRx3dUz60BtnYCnhtuyaTLKW2DtfLdbiWkIbVh6
tmaJxsNfmm1lUSptJ4gpi05fh07yzjurb9Mpd300Ug3qzbqOyU8b+1jH8qcaQGyr
CwLqZEJPquYUsv25NDs/PV8YFA1AMyBsItXkm7DmTpWzv8YQX2eM0SC0Yu5HIqht
jijdGBC+Q5ygMxb8hv3MG0GgA4jglJfukZdqHuYdRkksWhQARPSEw9dS5t7juDP0
bPsZ7EDIY4KosGVkQY67W4gDncl06nnbQOniZiUQkoOoxAd1N64qywWqcJpyZ4eE
GREHB2dGqsrm8OQu6HmB8Qjl013LX9gkvJ+A6Ij8NJwyf2PROq9LGdaH9SEJYAt3
wcWc2FT3eTklUejlFEknk2iYvF1TYXDxA9Fj0Axgam9sGYwllcHAlisyICb2qyhk
2fX4/CJbRRCKoqja0OdGSpXJ5kSuAjkVe5dsFXTBRfD9u6L1f4xijbekCt1gCjXY
uKpbWXwIpEPfw7J8ukJdBQm8lXxXJaY1LQIZsrC0o5+x//G/SINa7NT6u94pS6X1
Bj0v//uXLefeoy/M/V434BCBo1kFkO6kn4/17CfSArS+aJxx8hhKVAQSoDQbjOt2
KqXNx41cMPHalMnoNij6PCMPOgSCJE5LPh92lcPYZ2A6tnm4ssFgkDT1wM5U39SA
P7U6oT1lAXHYJi2+kV12lAnvGZ1QnVznzl2zNVBzEsF2l1+7hyh1BA/MXqARU1Om
il3hsOl/4oNJdgtC4eLYos1bv9VHngNNVERihCTIlSDE8v0vntlZAQJ1ap7O01Zh
sPXzIBAr+2g0NtcR6UVxKF+rAEprIW4JUhUAN/84N7x+DxVUXaST5u8VFKxYsM0E
ubpm+bFRk3JRFJtG9jMts2a1aeJ7W76PfhhPwkSag/ce3lmTJhbe1EHvwXCp/hCQ
dOhh6MIfxhZOU9BSe7A+RJ6+y1fqpXFY+ekLsMFi73tFRqxZH62txnGUM+XyHsCU
7fe6hRCpV3QHHU7Tz2BzYZUCo8sm92jLmf6nhhcZg37SfDB1mxkA1rE/Soe6eDtM
hYScQbk+5qfiC+g76TvMhoHesGwUk21uvzxXu1t//HVqnbwhv3LOpSbZW0Q2Voc4
N4pdi6M2cSdY/XrQ3hge59OC/n8EgHfEUAgOSR0tu8Tv7AuCb/amm9zsrL1mVgk9
/h3p75k2W21vVohwZz41Z7thdcGhMzXg77Y7rqh+9nEhRhzId/DyVn7ifF/V0+81
iUdNbF3KS07s3OWJJ58QnwCtvldn+so7xKqA6dlDui/ekfNIagQxbE6gZfqVEHWu
mkyxq7e0zaOHz/3H5Rwyv86jvc2Y2i0/gTv9d9efGfL/x4htPbxb/0IfqtanZoD0
wubmzdfO6CJEW5iTCsZgVJfiUZR/GUXgReoXuYbfvTf/w77pOMbM7IvV3KmNuaZk
29ybIb/0qxvqFBp8bWAnTQQENx+XGokkTogEnyW3uFB0ZKkLyTq5EBFEBlQmxofx
qJxaa6UFI4jUCaunojwXARrYIMA1YMYyUzxHuMPw7QeS8MNX00RnOBYITg+6oFKd
X9GJkTj8CbL6GccFK4J/GkHtVBb5Ve9ZP0FL5+XzuKOWBq06WF+XBjBwxVet0PVs
OZh06RG+P46R+gnDiuN1v6VgttdW6gMxdc5R84dow5L9LA3Y0xWECz06Jb7oXSqD
prkWOiWE4yQonY7X89Q2fiWeK9joRBomZVCf9+mtxn4EhBrfVcgrgIPmBC9cg/gV
MgBoe7p6kMgzGNq5vLKl9/FdqavvyM/zNsaxJjzJSRcp0i+RGcPgQ9zgqlULNIup
oki80FdEgSdCNLAtSFjHlAbnFBdhaQwZ6MBSprlDqyV7LpVYF7ctrDTANKubn52N
NPX7q9Em1sSCCTeO1CuytnwYJ2BKadBEsVd2peoqjJrErrDasjkf/1/UeNOxrXVk
kU7eFAgygFfegwVng2sw7yQq+USmnvuns5dO/nAy2kTTP36AT2Qd22Lxk0xCntFR
7mx9jPMNGVC8nNWnBlauPci0WdNYznDN0TRGWn10g41ejYFGE+un5TVOrSRZCVGJ
K8IMDnILhVM+ihZmfztBS8LiEZcNWPYX5Gsj8Dc6AihPsWrtHC7TGn0ggPaHU7WD
+VsWr7j3VpyGGI3EBnAtV+hUqLqc8ZrTAfMDIStwzu8s98f0OhLIhg6l5M1D9ZzL
P//Uu7h+rtcCbpw8ZbbGNQrF9SAZbGmPG3sUv26PXLYX6TCdaMt7Hk7RrxGarbSp
hcAkPH2HMvSMxh07c+VTEQeF9bDMk8W9D6HJ+zY6XqM3orIa3oEVDPTSVJaUe/Ja
+/EavO7uuQe7TK2dsG7VcnZKbtgPiHrlG4BLFGrR1Zs9N3Y1AfVrlwWKTz8PxN4I
5WC8kKiubsKtv0md3knFdiX3igJj+YOKbd8GqCBj0opux8RBRLjMOfjtGBjbf001
sd3xG8GFg3hDGZ922x4ufqfxO+JGQJWf4XWYf323kc4nQ2UOgho2p4HB//4Xmyqr
uUcPRrLddcaS19sIN1aRBSSHo0rGZPeX5GRutFPfMw8Zv7FJby5RDbvBFC49ZaQx
yH5mQgfnT4T/42kF++ZnGO/3L6Sq80PcYG+wqDqBfgTTsuJE6YtZ3ling/YWffG/
WUM8KdOYNpxOXuB1+SQYAzomZfwQYDT53MXf4wk77FRJ+d/6AELQiM+ypxNaHf2D
MTJhraBb2XeHho44rABxYlW4a/lSxLH8oCZ85Gd/3+dmn5pi2mPkml0NFyCDaKSD
4y82VOxDs1PrkBUsA3ljV5nn8sYfR84y9DUmTW1KnR9i926tSpwlq6B2oS/Q6AzM
jWWMdj+HYdrRaaBNdtQdrjd48ttLNco8Wzg27+KSi3LPD8LdzmSwpTytfrHHz5X5
+gtZUxt4Uo1n1wFCXPgbYn99lrd0uxrMoIl/FwPpXi7OOCuXgCBOJZ9Pt97zjfQj
xpxFtd5BtCSUUcIJxkbOlfS45CeK8DNRG3gEXxpx2pDOH0hQuZSrf2NsA9QDReL5
i7fvE+vxsvLqHwSp4y5f93XGyWqvHAaAboOU/sSEZVD1NSNbq0ve15AY+IwaJapb
sAjj+ZtCP0pPTv1YOMX0KYhCxgHeC8+DbyhyGYCU6UYJSsnTiiHQuw/XHxh4p6QI
9HarBrv/mJSSn6+U9NiS9OU6AuhQXFSUdQMaYmXUrc8+0Ysp8v2hI+ucEG45Pp3o
UNHtjTM3NPGyFhfjhYJJjlQTGzZTRukmtnJ5QE3U3E2Y8dyzs0w5CVMwlVRhU9ie
FbyQiz5R5QTCobDwYc7f37JyaXQjJzzuVsgZITMrgaaSfjBzWVu+Re/0fHYItDTH
QGwJ6G+BN6NsH0uVoN2XneNsdCY9b+ssbPwhON9ZehgsRQNWbRXw1caPW7zBAi0p
WtywDEOl11sv0d6S+gZtDqAKQc/+YH7Pl6AGBtueHgIJi4+RGMBVWHpy0IW88+cu
DWTrfdGoiOu98zpmH+fg4OgF+thdGAsQjKuZbn611Hwpbv2fihUcBWVxH5UJbF1F
ppusFrGkLK/vz/4jO4v4iXUsbs+VY7a0U3olGweZwb2xTppDMu7C+i4mGXZFt1mU
TbIi8DjY62fg+VrtVA8lUvWtG7M53BfvZ7IUY5Bm1okQed58T0vVQHKKV0b7Gv2F
2WwyFVWd5hy7+J5l39BMoI1X73IPv4Oynet1r9BimqpGUL84EfygTFvzKDLHYBc1
QZk0eYyn6htayfhDWSAFKCbNRubrzp0l28CRUEVuYELQvLOB2be2K+5yAGpOujhp
e2oY1wciRV48qgmHKKuMZJhJIhCcOwropB7hcw5La+STB0xF0XikQ0dpV7YRr+vT
Weog/4zKFFc/T4gCX18R8KNsqjJT4ftgwSDdHUFvmzzy3qigfiNReen0OVihL0fP
BdjGcm9eo/sb603ydV17BxZMKI2zCPk3f6hNubMNkMyqkANoQWnWEN8KWrT2iQVE
U7zDEPPGkf7nnhz4yx6KDIUnm05UtKk5p55xAplGBxggMtBg0S52JNmLUViD6Txp
ekuawHE2JNlcFQJm1TwdLSHMni0KzdGxuayanO10qb2lgul6pR7zqU1FQA7IDTwB
nfEUCxt1bcarxCev5x9ZhGo4a07nISg6RLPNsqGldyJNepJDhhCpTq+irEAuXvU7
jpsfQpLKvUKEor7c5MPTdrSeTSYSuqes8ZeQY5aZJ5ABW/Hel1Gj+b+vtsmwqhwJ
VtAl+Njedw4U+Tsm6qyKSyYZQRUrK4q4qzeZmMyzFTtq7+7Da8gWFLfupZHHmRgt
aiS9K5tS7ZNWog93cnG5GjZEjH7rmtWtJlakXcDRIartDJtX7Qzf0l9oXfP3y7Ip
w567jCdN3Ms7gCydCnHD+uvkd5T/Qfi8AWxWt/2UKWlSgZutOhEU43764cpajtP0
Kv2lt4Bd1j8RxeYUvPFZnI3N/W6CWfOteDHRvYKK6g34BKzoPv3O+AJtYIW3o5TG
/SzkPvQ6BqT2o/g5GkbkmvNeSN0n/1wIvCp5wv9BHh+5c3iRef1UZi3EQI/AMtab
GHul42+iEbRBWA3mRa3X5u4guysVpvEFCtJ/L5L09cOqslryoKRDrkj1rmcx+5cE
luQ3bPATnYg5BKa9L4hRrcgqQCrHXkM8yI1VC/z/ovPzK+khe72qm6MAsiRy4EVS
u3Bja9y/RzZgt8pcZtdTt73NCGsb1uMO7kQKS+DirC5HQ7a8ANoyX13SvjgzMuIj
KZBtX1EPZxcEAyw+5tdfnTZhfS6KHujZ2hsMMlO1oPgTwJu0REvdzNAyhmZfk8QC
8o22tmvp5bsNZLQ7eGBfUvh2JqqGCIcUf6wnNQghfq/SdN+A9A8SZytrRT4UGb+p
S7igHpMXNsEIGBPN1CDYoJAPu5GeVHnGdOIjcivjJKksFQ/JAQoGvlV+tJg1iFeD
5kaHRNli+grdG88WajnG0gx3XG+OVUCWccUi2P3Ny7Q46BoD+Nao38baP2DlTVoA
2pc8H+CT57WaBSKVn3DQFpGpY01GImSIc4wJQCYIixLfduBbSuoJTXNnftEiD88N
2gM2JpWFIrQNVSDYE5z9AWbzP9BY3wGDXg8SgtZ++IJ4c1Sh5/RNam/xmOb8lVhy
fWaK3MybAvKrqIz1DWEpxc6q1esylOHUC++z7ir9pPHhWg38cOprlYWjyyY4mYaV
veUrSVnoT8QmtNmB0qg0lwyxL3/a3jYuPHJEZ19CWjfvbN8/T4T/gixzgqBj2i4b
+YuoXp4AJEnUgBn4+pcBhAwVfswigNJ0xIy3DAKJskFHD6R2PGTS+BmYgKdBbHkW
n46VWaQpVaQ1Wk+YsmlpFFmdkGy8r6OLAJbwKiWLQ5e9gOn1v3fKCe4y3EDRWz4N
phEX6SruX/IA5xpteNHbTRibhFJNXYu9xED4R2wLvDHydhuIZLCdpS+cai7lP60o
oyDgY6rq0Usg/EirE3yPVwZh+SjDcx703sZhgpkjrKhNzlsJjcN2GKjVKZI5FswU
bTZQbht+oHzZK+JfbrJRJFzv/CgHCPigiV1Gf00P1PnQ6XFuQP+3cWiND6MqkKrC
xmN3WWId3g391Q7GA27Zb5gA/I+NTrVjYESDAO9S607gPtIh8SJIinYnM4Zq0B8F
jeBfgIrVK51jiss4DdjZCznWegooq51Jb5YOBwYSo5obOvfGSZ3OGh6sedfNoj1k
diKnQbrRpnll1pYcBod27HNWAG3ENJSP5gET3X+ZAbg6WZpAWoBESC73GHvYIhKw
q9baZWelNNY2wIpFf5h1nlqk0xDpT1yCnQQhwFuzTG9Fp47Htt2t5f0MJEzaMooQ
sRCRFjI1dkSGPCMkn9cfbFtzZHXJQvU8xo0sNysrrrLD/A4TJdhxUPV/8ZT/9fTK
vOoNPvSqoDMwQEuL85kSH6V++aO2PJA6VHOUIaAYuOERpDAXop/bJScSCYN62QHM
oHmb/z8oiXMYvevmSUM+FL37m8CTrwVjD4kjpsWLvBySq861uzyyqFoEqAscbPFh
M20WhpwHHFNMCJVC3GzuzvAt3EOJxC1Z2N9LYUnK1+UbD0gLeZnVt+bHdu6NLQ+W
GwtBgM1kpk343GGImBCGsufx1nAW2y2LJXhwe4sq8A50oi7YZcouhjRYJ8oYkXbZ
hZ7IdI/T3czvuxhGwij5gmoDWAPMKkNRXhPpkkhx3BjU0+6nxFDc5uhkrIac1fTW
CrhY4pVWxKSi35ULSaG/+gVwoRTg2crfXxVRqTY90KMiSDN7wbtIjKDqXWnGiEAl
rFhrYE5S0u2aFJTD1yNVeCdC3K6K+0dsQJaVL76QzQxfD3G7RCFW0nyCCytliS7L
5tvfw8sVRFLSSe0o8mfQKaL9ESA3qU1yCINW62w/fCKttEP9UxagoNEEoAOFwAUz
0fr2FUMlDOQFDTa14XeoM3e8mqc+dbE94BAtgUX+z3y5qD6NMyd+BrDCXM14ivEm
vmJKfuSZAUWiwOndMAc8AgngN16ULte/B2BuQUaraqvc/sdsDAP2xey1QbROhn/H
VNIynwisxBN2FDEti4+mc/1Jivs1Hc5J9vSE/2tR/xryd5XoG2RAZTkkevktXlvZ
hKxCYThieNtCR0MkrkbzfUh+GCqR4ZJ9g85efkHjs8BmtAdM8AQ1quJPeTnT30NH
MF0xzii9l3gZ1jTqGgYY/sQYB2D+M8yK38d6DRMGDxC0EzDcmIR8uDiQ0MyHVcKf
kq9fxf05D32D6ifArSh6mktn1yClIvUzx4NTJZH54Qp6U3FAGYKJ+2l7jPMxVQUf
CcbljT/yzVTaJ1Utas5jQznV6FKmIAC5K43zPWveaBtIcwGSdZAxmozycDuSXjCl
5NobxwymF297ZRHKfjjq7kELDRdjvf/tEmp9dQ01ZRgFfneFKacBJqlIf8O1VmJn
dPIMmpvU2m1Ii8qlBFgLr42eVdvAiFpLs9c0O9dg6l04LexUXTnHxYEYXhKbS+5E
dLlJRpUQKQjl2IUqp+thdp8FAvx9mvqQ0YakS4Rw0DxHlQJ7v1xmP85OAGF8WDUy
7NoF+t4rjDQrFprYoGfQgz4pHYXQdI2mlPJQn/mbCf4+acVyYTDmEGJCRmH4pkg2
vw2VJQfpFKeF2zw5nWTsAkpKxUuqnLF3psSOkPYhh/VUkL6Db4Dd7++8yeqY7YXf
ByEKX8WiFix2xsfjsPe0ran0INyZCbY7movmLqLKp1cjow2qokeQ0Bquyap/Bh+Y
Oaq0vzHCMUlWscw/MzuqK2V2wDKzl6pJkezGQjQyVAgwjcwKJEWFvL51strjT4Rw
19nws2MOHHXzoeuV5holfg+averp6ZkOzbvN6naHOJHA+h1O8kmM+f7RC5WwPqrk
mlRLephXE6Xy7IJkehQiYsgYx4/gUuL/IFogdA62ogbovrQzRMPqDDX9SfsCvKSx
fpKp2R7LmI1xpe4lYZvRAqVeDsbdixrjoL6dCYmSXnwWgHIcbo7IqBOJbqt68VFZ
d0uMp/Rx+IHarOmapbdnd3KzPbQzpCLi7CTAzf/yRprgMpbA9BA7cQqfto71gYL+
8sOIUXjF93goywEytTPv5z6Ky6paOCvlbK5EUN6ys/jOzheyRt+ZfGrIEL5zJDxI
RK9KiRbFY8Hp5PjbQmRD4+UBwydfW89CtnYHDsKfaPlboEWmCtBMVDZfxpNlLjji
5CVFvQCF+GlN/3+MXSAadBO9sgaPGSWrOZjO6UUC3S5kJsz0FhL2oLB8g3JY6yqQ
QMtjEweh7HXgRfec31KMbCNhJuYOhhhqe6cL07CfeX6YOumG8JkC8hW3KtNTxSNL
dOjp+HnqE69KdZpAIIDXRnYNBPrf/r1Hg7VVY+bG+9LvGWOq2Cm78TjoHqXVuGho
2FIlPLRBMg2Gn/IGQGJolGlu7h0smdD0T2v1xntID0sUiYtSGGS7TOXb20pqTEcL
xhviAqnKm4fX+S3CBCnZEo2pyOJ2d/ghtWZ6i2jqUYrABXNtyPA064kecdwAcGlm
OZEFoE+BAgUnuJSsXdhZfsi61Zjr8KzlOFtUWm1Ss9QYIY+c6uoMGNokMtlonaxe
6ihNY0s9DNvs4dTF3KhPTmuSiZex1lgTmIaLNjvOrFPup/jzwaq7nloFggH28Sey
tOh+qj9WTJBra7K0U8TFokEE7IKedgtAWRwRngh/yngDmY3imjznQW9dhePgteyo
UpIUAcfW4rS8jCF7Bf+jlRvFCYPAn53axLlRfnHmGQBMrMGbNAIAM2+NZInZnbMj
PMi0yIxQzvf53WglwKKS8u/hnHuGM7bZgDC2nyA/E1whA36c7YajY4DkEqGLKs08
Bq3ARwrQyVqiiUWafKYkKU9+dJdzJH8hwMaTfZYzxqLrcmCr/s7+1MBNDu/mRSxd
7MQM7Bv1cJ/FcmktYpgeSzWkXJXy73gxWHbQvltdx/Zcq8WffHrkaiIb3LZO7KZE
X1Nyfg5ynGeBJ8ItqYBUvKFGdIIKwrUO7vql+XyUmLXYRU3OPeyPbksvfuF6GNjZ
DXxbhUqIwUyNIJfEX4ooyHKf4UIrSu1HQFc6x+iDLiaBWxI+8/a8lV/u5GK0ycLh
5VG/TCgcCGTN6o33jFUtptNQF0OuG8oEHL+Uf9c+i5bVzmsGXb4RWP8+573pFSU9
sjdQbqsKTP7nQxoxh6xUCuxypWNihVF14ZZRqRKOn8UwVIcE8UuGsTjKe/21qyEt
rzDRGM0vqzCgG9Z9N3u7wOagN69zX4QsedTtTu+ooNtoke7IYJ2g1/EU9I2pccp9
N6w3EDUz3AW1lVLQXkiUjU3MHaNEqjI3TAayFTtanTyZXtvuCXpQ4O8XHw9TKk8H
DMTXDFCkr/DqojKiA900Wwm6G8eQp7vY4NRS2VQyliVb/UyA00RcY8GxhLJ3Koex
yhN2mJacrWJcluWH1udP3h/98zRPd0US9ZiY8uM5TFhSY7lnYQZpfyRyKvQLrnSc
DVnzP6KrZTQbae4oy3Lq/aMcDgidFlie1aYbFcGNoZt6TX0WHFxset+poGf1nHwy
hzSlwuiQMyZKOlz/qPLFN5x0Vq3DF8Y1+mVU8C+8izcnKoQwQqMMTGdLGNkFLv7f
+HHSdEIkoJGE3orsWRUNO9vDmaFuyPI8vwIvW1CrxBgPN5yNc+bKTKJgoXFv+0YP
8efnReXe6MwnFQ2AAEMk79Bj/lPXff1rihloIfVoXQxI+CYQE7xsotWX7vzthlDD
S6fYnriSBhTnDM+OogcN8KaPP2tOBorMfA00TtyUbahIH8KnpbigVNZhHBK2T8Ht
r+yZc8qMn1ikDM1bGUvNdW7fiAF5V77s0MvNGX9n/WNLZXO/7LXldq0kPm5mqUIm
i473fpjitcMAX6f2XSBmAenxc8Ac+s9d6yF9KVkDs0DfrVaNbDmlIEajojv9nDfi
rG9i4V65DVgI+1l3wqK3ptlnf6BzevpEjU3ONHm1LcihwD7ZGpfS6FOriDqC6YNI
2DqCZMG0ypXPZ0IrYvNEjjdwqRm4beVoYUa5ByuaZ3iJVSLyGz6X0w8x/8kXz1dS
hiocB8y5lG5OFZpestajwRgOxuwEna9hT3u1QYCoJ1U3mKq3QUy+Ir+e5YffE244
YiY9F2xt89YSP/hm/JnikuiTNUZArL52afT3ZzWiwaG4EyjeNLmzHdb1aVyD1wgl
urh9Aq+xOR9NvDjAAhXQLYcW/TgDyHhwOeeJRUnlAqO4J6Jdnlfc8lPcWtIovnWw
eEVQ5hJsHPTS8yrx/rzaRI25DQkyOMUqmNn1jUSrYrkquj3o7vMPTN8PnPPclWOS
l/qOVHgTMEM/6ptxkOtkNwqhptcK29PzNHQR2JN6lmLK37w41SoiQyABbu/wbHXw
t2mX380TIX23yK9WMDmB78XBaOdrRfy/YXzRLf3YHH/GNQYKirkISuKF6uAistFx
e0QSF0QCJR7/zaGu81qNwI5lIIs2KletsNqGsHbqRNdF1blp9j7MK6WR1UHxWgeO
AXpDfpZFOik4iH8C7ilBweAtGxSTVWK/PmB7HadMoC6+nqSdtdvu/QC4+IbZ+TYa
vfiQoexq4AawPuO3fR0in48Z20QwusWoVPlh/kNMnV355GfO42pXa0a3GC7VTrHJ
B6bIhO7YBdDRBWRbDo/rVmr3dkeQxVxJauWSoYwSkf1cbr3DfBAt3nxaXJQuoTgj
6UQ5c2GWxViuV28vesjn48GJjnsEmcF2feVMXLNEIyNLKYi+83cYcmY48WGfo2Wn
NctowDjJbvR8/1XUPTYYi82uXMtEyB+C5ZDHU/B6TrkZKTYAUyckojI5vmPjkprH
FYaF2PORR+z38uPvKvKkCY8bxwG+WhXqlocevmxaELFpGBVWvcgAppcPn9pyXgsu
WhPXV2WnpbZCtx3IQBs6osOkLObjs7OHDvq69o5rdszy3eiPtd0susz22pVOfGTr
5opvOUaNw9L2JwSk0wDWC6qjCFEHNNWqUvcL6larFNTzQVv1OWAehlmxxOL0nWK5
Xr5ojeqzutp2ORcZYFrkTxRwqzkXLrCc0Iei9P2O9+O8lsWYxEt24xr8RF2cIELw
9Njg/eD+EEwdVKqKFGnkZIdhZQJP5NMtKI2taDlUuG7U1pvIx8p7No6DeFM+qFwL
4ujXRJUcztWweomF4YOqgfyQDePdlyJov62z6wrVGioOUgua875fwdH44m1nK6qv
UO/XMRPB+mcYjKRMXqPH5Kqq26OsZ4wChGK3M/aOlFnEdAxt44DraMtvgZdG8X/F
eD3FBj5MNARCgLM8ayOVIfNBLsErMZQ1UZvXwctW9/OcSwC3MBEatVGOob8vqsQj
zPqLLGhuucBqbaBNLu4060DB3g6q/cMjRpzP2RAvJVJuP0nohTr6jcXh1ZRoe3xn
taT2WKLFBeVOplYoB+p8aCw1d3PBjrCKFV5xMZVW0BjzJb50Gql1bC2htPR+hx8T
Sayp/JbLvgItOMoUHKYiRCNMcKn2Roy9b1iHALTaN/rUJeIZRRe8gCt/lAGmnA5m
3FdAyE16gyGCHeBJ9w0m0DRWXLlwmGnh3mBnTkuf1nLIt01DWKiesCI2nxQ3Ar/X
pKprWZ2whuEmf4hUTEfEZ/Tl6PrTNJQbEVhxhmj6yIMIRIoN+4qkG4wT5KCqT5Fv
b+DbRBN1f79iItbNk55QmZ7xYZPprMqTuxwXs5JJ8/tTlSnviiFHO2EUxMa4Bv98
oCeLHM2O5EiWMHLO/PGuUE6bWwwtyZAP8dQegsxueL+hbcjEQgh+RVcGh4v6LUa8
Q7BjoDE9pkkanjEBDChbgks/LWyE3DKLP206ysUOSsFfCADOs6XS6f1M4Nru3XJF
dOhDGC68dgPAjEL0vdl0M4WsbeUZtUMUsx2yejAliOIku/VeEuo5hfccnkwbygd6
fOZtG4qEAYj3h0eQH3pAid34Schsn+3nQHO6X3KTJ+i+xiIfeogBfYbC4XTXXXb+
I7m6tA/tYuuAxiNHVeTkiXqocp3/xZNrXKc9gHiUrFszKfb8jmY+S+HPtUdSgurk
ZGsQdcxmm021bDXQN+xlmhGoeSG+DF0+93yplZLfOV+I+zeC9SATFzfCyg6ovT8y
W1TmYCt+bRmceSQ23MOa/y7YyIO68tNCXlAeRVOZ5juuEYw0XnMdwyUOiX4JTmLy
EOcoQ+jQLCq6dcoHZ1j0HmCmhnXImNs/TgWAiPFu1/JZBRHf9HLIg7AL55WdL3x8
y8co4sW3Mh0zhVjp9YVtP2hE5NjpZC+1ASZ3esPokkG3Y0fmS3zENXb359SwQid8
xi25lNz7vqqBfH4M+36UgyVcOnw26qCMMZ/aZnjRHS0kbsRMljMxJyL8jv/96tO7
//8dk5pDOk9XYQ7IG6qBLlh7y0zxnWmV48QkqwlC1fHIEXc5WNx/3rNfK75Ligi3
2IQb1aLFS+hd5x8pvgJlnyMh+l3yoIyokHsYLDjUBXAVD06uHod2mUnIvvL1HX4h
5QYKnqiHyuVGydP40URV841t3swEzal27BmRR7IK9+ubFW95LG6jp6f2LX/EB0N1
1Oc6ji/g2vDzau6oJ7SSQ50QdZKnGFIULPMEnr/tA7hj64bu3UKFmCgcPdZshUyN
KQZ/tpg4wVUxA1T7F4DdkxLdlfe5WB4MN4BGOQb1a3y4i6mQOGT2G/ql4NZDR8oi
4nTH6jKzepNStjJGQ815TxzrB8RLtgj+zYL5bccbS8PKfYkgUWT0c2CnvoTgn4CP
vaZb7/RWDhUjhYFcrL7VLyIUzraL2kK5gvczaSNEFbtVP90BMr2ZcV2VrMzZBxyf
gvFYE5dI3qNBZC/Gnh4u6uKiqzgR2gxpJWRZ9P0uyJefBQXG6SQeAj1xWsMI8GYt
Vs29twxYEJrBq0N/IYK8AoYsYWRNyiP0m+rcw+Y5l+Q54Zsr5PV4mkr32JadKKx+
TIbgH6FE/VgGE+9s0RWUPuf/AD7jFD9oAXTpbvW+24HmeRVeBdMyBgGjPgnLg5Ry
DOkEjgPCsrt4jGPN9TvTLmqMLp5OhH1FeuycrVf7tJOrrcb09DoFlxyLVJEyxlw+
s8eLBTv1A45rENnclcHtyg==
`pragma protect end_protected
