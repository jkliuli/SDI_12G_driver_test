	component sdi_tx_sys is
		port (
			tx_core_rst_in_reset_reset                  : in  std_logic                      := 'X';             -- reset
			tx_phy_tx_cal_busy_tx_cal_busy              : out std_logic_vector(0 downto 0);                      -- tx_cal_busy
			tx_phy_tx_serial_clk0_clk                   : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- clk
			tx_phy_tx_serial_data_tx_serial_data        : out std_logic_vector(0 downto 0);                      -- tx_serial_data
			tx_phy_tx_clkout_clk                        : out std_logic_vector(0 downto 0);                      -- clk
			tx_phy_tx_parallel_data_tx_parallel_data    : in  std_logic_vector(127 downto 0) := (others => 'X'); -- tx_parallel_data
			tx_phy_tx_control_tx_control                : in  std_logic_vector(17 downto 0)  := (others => 'X'); -- tx_control
			tx_phy_tx_enh_data_valid_tx_enh_data_valid  : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- tx_enh_data_valid
			tx_phy_reset_in_reset_reset                 : in  std_logic                      := 'X';             -- reset
			tx_phy_rst_ctrl_pll_powerdown_pll_powerdown : out std_logic_vector(0 downto 0);                      -- pll_powerdown
			tx_phy_rst_ctrl_tx_ready_tx_ready           : out std_logic_vector(0 downto 0);                      -- tx_ready
			tx_phy_rst_ctrl_pll_locked_pll_locked       : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- pll_locked
			tx_phy_rst_ctrl_pll_select_pll_select       : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- pll_select
			tx_phy_rst_ctrl_tx_cal_busy_tx_cal_busy     : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- tx_cal_busy
			tx_phy_rst_ctrl_clk_in_clk_clk              : in  std_logic                      := 'X';             -- clk
			tx_sdi_tx_datain_valid_export               : in  std_logic                      := 'X';             -- export
			tx_sdi_tx_trs_export                        : in  std_logic                      := 'X';             -- export
			tx_sdi_tx_std_export                        : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- export
			tx_sdi_tx_enable_ln_export                  : in  std_logic                      := 'X';             -- export
			tx_sdi_tx_enable_crc_export                 : in  std_logic                      := 'X';             -- export
			tx_sdi_tx_datain_export                     : in  std_logic_vector(79 downto 0)  := (others => 'X'); -- export
			tx_sdi_tx_ln_export                         : in  std_logic_vector(43 downto 0)  := (others => 'X'); -- export
			tx_sdi_tx_ln_b_export                       : in  std_logic_vector(43 downto 0)  := (others => 'X'); -- export
			tx_sdi_tx_dataout_valid_export              : out std_logic;                                         -- export
			tx_sdi_tx_dataout_tx_parallel_data          : out std_logic_vector(79 downto 0);                     -- tx_parallel_data
			tx_sdi_clkout_out_clk_clk                   : out std_logic                                          -- clk
		);
	end component sdi_tx_sys;

	u0 : component sdi_tx_sys
		port map (
			tx_core_rst_in_reset_reset                  => CONNECTED_TO_tx_core_rst_in_reset_reset,                  --          tx_core_rst_in_reset.reset
			tx_phy_tx_cal_busy_tx_cal_busy              => CONNECTED_TO_tx_phy_tx_cal_busy_tx_cal_busy,              --            tx_phy_tx_cal_busy.tx_cal_busy
			tx_phy_tx_serial_clk0_clk                   => CONNECTED_TO_tx_phy_tx_serial_clk0_clk,                   --         tx_phy_tx_serial_clk0.clk
			tx_phy_tx_serial_data_tx_serial_data        => CONNECTED_TO_tx_phy_tx_serial_data_tx_serial_data,        --         tx_phy_tx_serial_data.tx_serial_data
			tx_phy_tx_clkout_clk                        => CONNECTED_TO_tx_phy_tx_clkout_clk,                        --              tx_phy_tx_clkout.clk
			tx_phy_tx_parallel_data_tx_parallel_data    => CONNECTED_TO_tx_phy_tx_parallel_data_tx_parallel_data,    --       tx_phy_tx_parallel_data.tx_parallel_data
			tx_phy_tx_control_tx_control                => CONNECTED_TO_tx_phy_tx_control_tx_control,                --             tx_phy_tx_control.tx_control
			tx_phy_tx_enh_data_valid_tx_enh_data_valid  => CONNECTED_TO_tx_phy_tx_enh_data_valid_tx_enh_data_valid,  --      tx_phy_tx_enh_data_valid.tx_enh_data_valid
			tx_phy_reset_in_reset_reset                 => CONNECTED_TO_tx_phy_reset_in_reset_reset,                 --         tx_phy_reset_in_reset.reset
			tx_phy_rst_ctrl_pll_powerdown_pll_powerdown => CONNECTED_TO_tx_phy_rst_ctrl_pll_powerdown_pll_powerdown, -- tx_phy_rst_ctrl_pll_powerdown.pll_powerdown
			tx_phy_rst_ctrl_tx_ready_tx_ready           => CONNECTED_TO_tx_phy_rst_ctrl_tx_ready_tx_ready,           --      tx_phy_rst_ctrl_tx_ready.tx_ready
			tx_phy_rst_ctrl_pll_locked_pll_locked       => CONNECTED_TO_tx_phy_rst_ctrl_pll_locked_pll_locked,       --    tx_phy_rst_ctrl_pll_locked.pll_locked
			tx_phy_rst_ctrl_pll_select_pll_select       => CONNECTED_TO_tx_phy_rst_ctrl_pll_select_pll_select,       --    tx_phy_rst_ctrl_pll_select.pll_select
			tx_phy_rst_ctrl_tx_cal_busy_tx_cal_busy     => CONNECTED_TO_tx_phy_rst_ctrl_tx_cal_busy_tx_cal_busy,     --   tx_phy_rst_ctrl_tx_cal_busy.tx_cal_busy
			tx_phy_rst_ctrl_clk_in_clk_clk              => CONNECTED_TO_tx_phy_rst_ctrl_clk_in_clk_clk,              --    tx_phy_rst_ctrl_clk_in_clk.clk
			tx_sdi_tx_datain_valid_export               => CONNECTED_TO_tx_sdi_tx_datain_valid_export,               --        tx_sdi_tx_datain_valid.export
			tx_sdi_tx_trs_export                        => CONNECTED_TO_tx_sdi_tx_trs_export,                        --                 tx_sdi_tx_trs.export
			tx_sdi_tx_std_export                        => CONNECTED_TO_tx_sdi_tx_std_export,                        --                 tx_sdi_tx_std.export
			tx_sdi_tx_enable_ln_export                  => CONNECTED_TO_tx_sdi_tx_enable_ln_export,                  --           tx_sdi_tx_enable_ln.export
			tx_sdi_tx_enable_crc_export                 => CONNECTED_TO_tx_sdi_tx_enable_crc_export,                 --          tx_sdi_tx_enable_crc.export
			tx_sdi_tx_datain_export                     => CONNECTED_TO_tx_sdi_tx_datain_export,                     --              tx_sdi_tx_datain.export
			tx_sdi_tx_ln_export                         => CONNECTED_TO_tx_sdi_tx_ln_export,                         --                  tx_sdi_tx_ln.export
			tx_sdi_tx_ln_b_export                       => CONNECTED_TO_tx_sdi_tx_ln_b_export,                       --                tx_sdi_tx_ln_b.export
			tx_sdi_tx_dataout_valid_export              => CONNECTED_TO_tx_sdi_tx_dataout_valid_export,              --       tx_sdi_tx_dataout_valid.export
			tx_sdi_tx_dataout_tx_parallel_data          => CONNECTED_TO_tx_sdi_tx_dataout_tx_parallel_data,          --             tx_sdi_tx_dataout.tx_parallel_data
			tx_sdi_clkout_out_clk_clk                   => CONNECTED_TO_tx_sdi_clkout_out_clk_clk                    --         tx_sdi_clkout_out_clk.clk
		);

