// clk_io.v

// Generated using ACDS version 22.2 94

`timescale 1 ps / 1 ps
module clk_io (
		input  wire  inclk,  //  inclk.clk
		output wire  outclk  // outclk.clk
	);

	clk_io_altclkctrl_2000_dpnsueq altclkctrl_0 (
		.inclk  (inclk),  //   input,  width = 1,  inclk.clk
		.outclk (outclk)  //  output,  width = 1, outclk.clk
	);

endmodule
