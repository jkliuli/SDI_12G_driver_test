`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
cZwiy5iObAHIHTxlwNt7LMsIRFZZb6RDfmT/KSExaPjlCn56NrSFaQRuQEzoxbIS
k9HomN8qypuT1FrPQRUk7+AjZAdmL6KkwdSBAt/nOCs4bA//g184M13qOSCQ9Q50
4MUlNbUu2qNkrz/SSL6SyWxPrm34gpjc6D9sBtMSUis=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 70496), data_block
/Ca5zRkhsTugtEFMjzL2ACAsUNXUL6pMcmeifw0gk8fxtxo9dybMkc2aoUs33rRu
zKqlmFkQooBymZ+6JAB5pBgIm10F1T84scZrdZ8loAoTDZ/KIWz6heigpsBAIaBm
Py3XZ5g2gyXWLcQJNR9kv4XmQSc7L670HKkXzpCN2Uy0NdNsHKGjdbP/jeIQuwSl
6/tvsWQg3E94vrtRfvV2AHIaMLtXmkRaQv1M8bIfWYAEmyQ5xZqAPj9bImDqndkz
1qSSSaIRRHNSABTlof8t+9NNtGStN5jlX2LSPqNjMo+dbrFIjPtVd0UGnxhsbiUP
+kufWrs8WCTTpQbOPWLwiCpE9TSOrIFZeIdsCb2nLL9Wzy+v/eY+NuVT+Iifo8KP
tGXYsk9uhEaEeiTsoWqrijtV/vN5h8yWD2NX9lx2eakh4QUYYnTFjpN09DMlg/u7
+QrzkWPd/Zc7zGlYMWW0WSW8b8ZjA4i41kui6rsiQTAxn1YbGGzHcqRA4tICnOh9
GdG3nIGpaDI6qeq5w+hTTrZh2uYc29+HPCmrkPaSx6gdGb8LEsqvTR7MV6qmsLGT
CBgKjUE7vAc6Yu70XuuKD3/OA3Dxm6meofABzsRNhw12+6AWWyHSzzIoM6pqEmsM
EHwYLI+7J1EoW22NJmHtFMqWh+F9NlcXAUIN6CPFnzs297m8spPpJYUgLC/eEErr
BHSYoS/MPUGs6NZHtSQKIEIzX6WdE7uNHTNtMjC+B0OfoFFEEyzJOAJYMkNFUS+y
21QNLTomWLf7xVveDbJP4MPSrxPLefyuO+sxxv4jEgxYTsF3fBuIrR7SFZgnvSRA
yTmK57KXVVHS1wkzyJFcX0u879R0vBoeZBBaJKZcTMGdO1G51dLeU0wjJuazVC5j
QwMhJpHilqOjraqYSzh2aNrUJGXFP3tsuY7butknQhPcCiyMgRhik5k9nvI5Msdl
vbdEbQW2Bb0FRsXiDoSZ7ohwrr1KinVc84a44o4pCrmaK65AGE2q0dmkQH7jhzOO
vt8LR822x1bnG2xc19YtWdvowv0gDlMHgcF7yV1eR7DPaRlm8Gc7O7wKd9MeGhnX
QRkbbLGIsdsegxihQm81IFjdvX1/CcKb5Y66RTxHEsVeCInLn1c4t44RraMCMTo3
AN8SfqglrUHnfFBTYPAGF99ewlDYbNLO7RA0Wz600IeRHKrOs2JihKMdP1UKZbIZ
KPYaFaaBciWf2+b247xWWyZ0a7GmK8eaF7z1t192/FCpLQx57BCLFdDDNjJ9I04U
qsm9nQzy7Z5FClnfh5FYEKTyCVoh5WULwFL4/Rqe/WJM7thREXWH/cV99U6U459L
aqiFt0ZMuzvWbyNfAEZPdIc97Wp9cjtyUEXb7W8U2EY1bcCD4/+do8JVEDmqT+N9
NCEcdQg6YFcRKtueAZa5xX2mQSoRr/ePN3AAQ8OJlYBkKXVUDoSoCrRSpXI13TGA
H4ZvJUrXchd4fdabnepk9Lw/fotcDUsJ/7Thb6w9MHt3d8+WjlYLexFiXsBZqubT
hmAqOVuo2E+/Hpl5OrGW5EQ5tGiX2JQKAXgV196QgrWKiY2pP3FOb0poneAyQvuG
38bmvOAqQUkf80Lt3k/ZmCMfXHyECvui2yT17zpQ+kmL3zpIsyo5XOI+6Ncjhf7x
48bfimt7JT3B39WQqVMHWcvslRopFZ0Qp2DSp+Dw9lfQhEUhDvd0RtJrWfCHd3+N
wozOTRrPZAi1DlvHki+gwiGa7i51j1dWWYywZorZunjHzd+k6QK1IgsGts6u1sdD
T8MhPtOhWeILmKH4GXrhxtRtPZlaDjFZvUqw3bk7vaHz3nsHWV0f2ppTDZhCr8Bg
AJydf+gbvJb8ql051WIlcGkajErd+qpnwTU02kjuT362x1RGPqbjfDAH5zo/lsho
lq/cxBeAKbo5/Ilq3o9/vMiXMJUjIjdwN4P48KcIMWYP4eul1UKS5TYBsL2Jaou+
11C0m+x4Wz6sg90Xg//MR3SyVHH9JaZKiVMAtl7tph6tvVSJ7v+Ey6WJXnzitWsV
1NhJ1M0cpxIgiOWELAxL4315ulyyaYQ+33v3+RNoMtxmDEvKYOZ45clpUxIgqQTQ
ofYqkZHPC6Mv+zdEEpGXmzZg1Pw932qpTvw3XiP1AqzJRJJttVbN+sdooEimlB68
ftpYeCYRm/cx4cQ4H8tKS/XPsQqtE16RG1DnbAZbenFxA32ITCo6f9OGMbipLB4U
Ddb7iOmU9OATnqSKAnPRc7cSIrrd69CF7mcOttVN7p3flqTURsJUi/nlvGPiQGUJ
4ZM462WenUYz67ZU08y0o33Acm/9pFU3MsCilVlnnvQ4sqteN7B6FSgrG5hXeYYE
fbGXqxL2KhbfeIij9M17P08Hw/upIxgBJ7sNzfUkCOeLQAlcX02MQ1ql6dVJhseH
HemqtzMQ+8cLAgevKq4k6wxzFyE9IG7ETgIZGtgq8DkvOk/ikrFCPrw7ggL0pdL8
mjQzjaTkY69+QpRvTRGkkTWuprf7dWHihLnW99ymX46RIXjb+46fedIV/6U2Ra3U
Kbwwx8p+GCegh+pWAsq7aMmZumwgHqEhnPiZ3XSUur5qpRnkGzLSFkptaQw00FSp
2U/uM26PykDWW1bfMMI1S64Gy/hVzcYAdYUlYCpVfgIXK9TBvnjS0bChhm3qYPlI
MxepgAZzo0rPvVDNeti2Xg1WOMX1iemltKVdqvy6r4HYfsG97+Kg1MOoPOVzTsE+
Y7lQfQ3mqkKAFp57YaE7Y9ZGeRyGWBIR/CUENyDRKVEDLHi8RoyvEcfE+GEKq8SM
Ia536Ymo7KljHxCCkP0yKzO8YHDM6csd10rcX1+UpaaBq01Kp11YdE4UmpaJYyMw
xRzgL7Mos5LRm01ojWyAYgjm1St5JsDmuSdM9zbEfsR2niwE0PoreKq0Lsqm46tQ
5r0g0vsxPXNco77bUmJFqLohgEdznSwqtzmdALSq82xi+xMF/OHs5ni+NfBhJ0Kx
HvRm4djHhzCDDNXVEyAn6oKWQat/3GLBZhqgOrG8LFlWkHS076t5aS/rRfkqU6th
E26sn0PRH41uEZT6e2v0pL4Hm1aoETAWGXkA2t7wZTQHcNf1sPufNGaNBZtSYNXm
nbhDF9c8XWnW7lX7wAt7SMMBzERGzhO5OOcz0lFYO/lM/c/hurm8oXosqHC6mb3O
U8cBfGE6fMPMpNyoZu6asPpQWCIOV9LwmNyEwvTEWmOtaLOZtMOFvr9lJNkHuQ8P
x7nAmbvg1TuoMSAokQ8uRCrXwS11EbK7n8d824tUjWsLAILz2TLJMCSYiOVw+N7V
JBDQK/q71+73oP55We8sIoyQ2XrHqJCfZvOeMByqFwM2HduGZFDMdsloxspEhwxf
G6XczDci83B5V+ODKq7tMY6SNcBlHm7HUEI7bfifuJD4EyuW+Wr/SbaW97sLWIVx
4v/Sj0bPTPYp1whmmik3PPz+6RANzHfPkMGTNaVw+jXwS3OtyIrPnoIcZ3FXAF1F
a1rGzWEbNpVJMm/k9HUcUOkRsPEcULC4zCS3UJT76zd0Gu0C5V6bzSp53O+FbfDV
0Ju4etMTKaXiMg5kixPjcPPvfknZ4gOSXyd0AAbYIouKmHV+fKzn2l0L6xVYOD20
Gy+7+6cxrlF/D9W0nq9Dq/f9Y0oHBODiN8dMV8/EEDVS/KaStqiP7VpXDq2Uw9Sf
BV1cgjsZ9xzAgCyYEatL1nSCusulKVb1SwWQxn0UzP+D/ZsTBqSqP6z9Tu3FHpeR
QzJzuqe4RaK6aTuIbbDRK5DC0jL2eyrTTWg7obKn5n9VIf/YgvUEj9iokeX+axkH
0xxXDHgWhe/spw41Uxvs5wu6vq5xjxrzk4WnzoNq1QaMA8bqPL7grFpYCqXzx7dq
zzreU0TQPjH55/eN20WdybQlOx72iQxWSAE1OWXfDiKNokqLF5DooLiswomTWTDk
kd9yTdyhCttbLINe+oWzvX2KzrC8f8HM84W5iKIRbPDYAc1VitKauxJYRe9vpvZg
0Z1x50jx746PcMTOJb2UoC/93tbzp/y+PrKK7duA1g4ZAWlnwZE2d+FyfEetw4l1
u2NQw72edGUD1CDWb8HgP6OZBQwlOgs0lDYyC1kgXAlswPh8jY02AJaE/7WbMzkZ
P0eJ5CRuPdFVAmveH2wNL/gbJve/ebNy2/QlOQhfx0pMVMMi5PImpWbNUgHc6VzD
pHpXq5boowJiH/R/fhdenJ0f+O8rWUbpudupcEoBqdyV+GH0BRD9QbipUa7JabOA
SHwVwa5y/HZOGNx18eblLQ0U2eoitd1qCnu7lFGA5ls8iW9m1K3slOyR6+We7ZBJ
SddbTuvpXbAnmVO4lX58uDf86GWnom3VyEC7yhm3nIiBzN3qchp1IuDnShQEDqK8
I+YMBXz3/xqYUgAv3IVwPfhugaxaFOJeKqHqT0HtnVhwbi6w7twPznNHUSBN/v1s
sCqKdRXDa5pLlIZh405JNs6w9bqMO09ocT2VlcDfKLqNV76/lEz66jZ7DLPxrhPB
DN7ok0DoOnFug1T6mhrPJ3UGxRyZzrcvHuL0eGoA5T2GoPQpaIBVprF2huS8k9sa
fgAG+nAty7kW8q3ucUx4gyQOPNVmCkj65rhC6Oy3dURcIrkmdRDksh6u4I4Wdxdq
NRw/A77hEUv0zRklDJ35pUDn9hiBwAjtjhINL27OPuKJsEIcM/f5V9081Mt+45SE
jZTQoUAAN+7TQM+KFZCnJWz5gVcRXEprnMSnOT1GLLquiIk1axUmTPm/Km66n7OV
bmzjqFujFwiZyQ5OifNgFFRcszOPth2GMtaDyD7lZna/K9lsvrkJSlLxK0N6pc/U
FZfUmwBTYfghSnxpX5m1QqkAHdqs4kPN0qOBU7N7A3jVTw4isKDxmrfGLDYq2brc
/3wU0kj9cevGeV5JaY+YVhEMLncH9ovKiLvgm+3WionlatI/ZFCm9HneoQLZ2VNP
mG+P2IpdAroLKAqVtVWa0Qrh3v4QJ9UGXpH/mAGGN/IVAA+HB9vLao2mEBPCm4YF
OycrcfuPmw5u5tPxWdSTCUWXaeNnkmx0snVRaJ74aNP5ioEzIEs4y/2kiMjOD3hr
E9Q1GistjTLqqfxU8RJ+cxFPjlQkMP2ZiHb/wQxUb8K1LLjp0fkF9aC82o7OSBVD
INoW9w3h1mc+B/hJVWNxczHUHz7Q3x0it9c+g67Jbi80b5OJi8Li1TASE3Jx76cn
psZHc8doYgR1X/Xux37PS5Vyi1XpuvNyLLwQNqeBmJUtci5bUgGTklJow3jxqkH+
UC/Woyt6pzeOyFTCNEBmueBQIWBWzdPgjE61J9K9aAOSw56/4y7GMRu1Q0DBs5zw
CJrjHydTMbzHNoAx1wcwu0UUQKo/kj6f0+EFAiWehqwtE5WOpwaiZL+JEZXAA3g0
XnZQkiNhzWTq+K1lUU3It4R0+hE+sKckLUsnhyxsPfdp6EA0NP72bVXZX7peXpdH
b6Pd9O4TdHcRekELnIpi0flRLL/DTPX57nU4z0GwsKGbAsJvEUhE3oLC1MLvtYUo
lJEM5psq7869R/7DVEgzjdoK5rvgnUhdQDcoM3eXYrfnszfDMrVjiT/UGS8U4bdW
DJSf//fYA2f0XuGAQAjjgdf7h6WfXwpOVSg3210vmo7J0L21M2wbAZ/XPDplF455
phQhAmQmhm5nANTHWChqqLLVdyMTBPFnltfOV0volMdG99z953aPdkpjZzSAnVE4
/8dpxBYKXoN+xIaSpn49smlKjTYcIdLUwGMCXQ5eW6hehi4/2pTC5qb7ga6o0R1m
T9WCIidfnKqchcrrMi3PW/RgvZNIJufPYz3q4lnwZUJ7MTJxiyXqDmGZtq9T4ynX
SdgsAQG6fPva60lX3nNbrVsqgQEulvDYar7pqW9Oj9do70KVIL5tZ0dP0sNfzioL
aHk1UfK80jyQIQEi75C+lkF01zCFNIilHPs+PBNl20wL/PD5hbhHZvEMpuTboNVv
ivEbKpVgKmrcVCryPfOJSSEs1t9NjkwuZMvKNbCi46XGXk6Jfbg6e6tv0JLTcCv+
aD1D3VPc2LafQrirkJf+04X+TBzWBIucnQTyCGNZ/eNtRiskGBNKaWZ4+Z45SFj0
X1yz2TLgOkGAhZwYA+rb5a8Fdw55E5tLHklJ9rBnX+X8IP7XLrgmTCxcmWE+ziS+
UPiqvVDvUq2EoQgma4OvL8R9ktfz3Vrf5R+89b/RE/1TU3Aiel4WoOM//DFqHB5f
ykFCFuJhoTJCCuGTwSpqdJOKbSUDKuJ4IN91oGD/iuy1xYfWf6IaHZdG0SHYXOwF
OVrSE/XWzuVXjsrx0I10ZUDIPI5ujsOC6HeJSJMwwxbRGuvmVnFpltVUK8WU4wAX
2mpnJJgc3wTZNJOScEynxLpRIW9wqA4JIUF2CLpZQcbApwbZ6i3B1Htkc6gzg1S7
tHINIsf9jcmKi3t1q4X2F4na6E8sLL0yppHEc/PkIEf5/id81h+oNP3WnoJ52Vdy
yFa2cG7etfD15fgMO/AYlzz2JkZMrQmEXcDJ8L+fORmoyayc5FZn3dWDR3M2Agtw
rSV+3uOHcCYTkMfqUq7osaxbQx/+hs6HqDP64xnh+xftOX+A6IcP4H3dU5enm7CS
XOoBfLIR9YYn1VzSxQtJZKx5oTZrkfbvZV/nyYYRZFz0nzJjmboRP2J3WPlWnev6
BmoWcRddThI79cDvwPC9zsh41k3YblmCd43/3BTOLgBbfTRYCcxExGU0JM1H6uIL
D3XWVtkk8Ua3TmcPG8TWeoL1KVHcEizjwTN1g8irkQa0wHB4E21gfdiWFfOel4F3
Z5cJfm11MLvBc1YXCh4GZfow+Db+VxoIiPPTE7v26KrLqrW0Xde+GRr9b72F/YYt
0CKBbQf0xLzkZE/kayuttIneB2wJjFMl7r54mts+Yua+wjNYJb7XhbM1vUILj9Bu
0cryUGwJ4DkghlXj8Ji0oEjshwVoMVdHx3AtVaw2tEHxznCKeqpzcVHCIrOLQ/f+
vgFtC/a8gKEYbjAizikJBW09eQpZ/CrL3E9ar4rA9E7N0EA8Vhz/muPpCMXK0R4z
KXI+COBqhxLIsGm0n8lkxWPjUxagplOeoKZudDrn7GqWG9Lbug1GdWQk91bDvbd0
xv6dOWEyYOV6lt+2LGQgCSkZQb7ecJT2ZpD10rh4byOXyxKodM4iJMUuhbU09A4U
NcmmgEMAdUrYawhOmzco9sR9WSDrxggXSjcEZmwq14fFScOtjnokVMsDe4DvWdJO
mjCuV0bbsIcUS4nbzmUQVerDSnzfg3yitVqvueOv7zSHEcwUc2+439+STX3Yctc+
wDj+N53XuwcbEwihai9x245uHwpQujxQgCd7Kv2I+qJPjbyru40M7kLNe7CFhLQB
p04ZHUXf+dWmAwRd2BZrHyF7YLeebzxuX0fiSdJgK8tUD7CB0qLYbN07Yk5wQX8V
VvHU66o/3rRqFwwnmrrkoO6oF2nI5Krwse6SwEo0n2GPfGyk5hYsfFFpmbsnFTAm
AESu0Sng/6QYAtcuV4QHiIfDLgdo6hnp0sZb7NgQZ04zKYCSEurPPWVye8p7o8wO
Vn9gvnHx7XrWAuORaSc6XPDqfuvYsdl7rfIKIIUYf6mkrEgX8gdoOoBeq6RbrFQQ
fhHR4EXfHk1LnBkAKXce1PK36NdQstmjn24c1Ic4AJLRDbgPxvucZVTYed+pGfxY
Go0klIavbFqQUaDo+mnrZohg67eR+NlPdrviOny7NQH6H9aPFjf9Am5vF8HRt2+C
lQlQwj/hFl2Ydusv5/Z3l93WAXZqnwYXvsyCy2n4jlzatirBuzniQ1SbYYzLCMBc
DPCUK1NpIBYkwdTyl2xa4ep1mzPooCZoL/iepHhsWASYJrnqbw4YxNdOxZFl32Vx
rQQBz0LjboksWNbQ+UBJAvG0ur+jSLrA8IUk6SsQwlfcynBRK0UiSBt5H0V+qtfy
CvlMRI8+D5mw718Fh0d5Gl3raprE6+LNN78bysxtibWtnXMOuLKSuaqzwU4FL5cl
VsiI+WhqKyr/shU8PCU+DZAI8GXZnmiy3m0U0dP50YOXNKzCQiB9H+MTMIeCT2EX
DT9KPrEznrCkiuOOuT67/cCVVEE/Zc9yxPIB9z7zATw4lApH7N51itnlE5OK1zSl
AR8tvlDNby6IiyER4KzafbXT0a8GvZbVA3FMD97WC8hA2CrqJkaa71tdYGWnYdwe
enzgbBferssIuILvTAQeUYfiFBUWn6z/8/RDEq1Mf5kLByP7seQK6izdw8Q9WWuy
7veFbhnSaec+Z5uBXB1FFMztgy5FAvB2WyN1MmhHerDZVyMFX8/Ur4Yo3dkNwG9h
3/BTC2Ar3RgGx849TeoOszil9/NEwwqkFzKOg8U3NMC82ba/J663nrfWfEXQS+sO
xBtsbauHWXB4iLkyNHcbohxxGAfu3zWoTBAaZWuNn6L43MovbHHNq2n128HdeIEa
HYFFqNZkx0HOVh85ZlPSp3LuRwDwjh7ThbaFUU7EMWx7oYlyaiOvHMd/h9ItWmva
BE7pgachoiAfFjj5Q7Hchhm8mBpxAI/rnPq+VwoWY0Aem36+JynBpCXUP737A0eC
RMOijA3UywqT4LvMLsgBeK7Eaz6j5f2l260TipM7wdaRBdy1uYpSwYwXHeoyjFa4
Cmnx8uCiYfPIM9sY2b+nyUs0MsHjdIH2H0w5hGWX+javORrT/QWgAgwMlvv+1FMb
h0+qDVrDVKNMXzmX7AZ3RCzRlWeNazlFrmBc6CygWHo6+AHfAdQdZsofGkxMYEiP
FkMK5+3dTN9nj3giWeUpy3rBsUHlWO2O3O6ttuUyYFj/rlYkpZefpNM+jNITlxhM
AiohkpX4kUuFXFGxpMAarccNg/shsemxECfxHGTmNftNZalgrg9sHbpZlblLHVdH
FvD44huAIdXv2w3VkiIaaSDuUUw8OITb99BaNXanA8YIE0AQ5F2EJx4lLRgrv8Zl
5vwQhHCX4MwUvhEXCnFXIpAkXOUBoXv8K+dowI5OseIusO9aP4pGNDr8r00G52lU
b9iyhO7tGsP5umRAUco2Le75at0dcBiXCyyxcyu/OZHMIBrCGrU4+GMw8lax8WaG
cQS/pIng5t6Vx+ulTEWsBxMSpSQrGm91JFWKLy564TNRtaROq1v3ptkZGY5FTBZM
lMtHCIOQZ6IykYvXhS1ixSA9BbXDh6iUhydDZuPxJwCSL6OiPeKWa6ODwDSYUk+0
9EkhbOCQQC/4X+apk1VzmWY9qLDv66EAFUMCiuSsUnZK+AjKH33frS2JUnqu7OLx
53eljYJf0DJBSkTw7q8jQyN2xbaT4t7dQjN7+kTAkARFu8Ey23r7258gBcjlHDXG
Df8HcIlIiUaHXK4149j4cUNYmyOd+XHPHA0XaHQl3u20QRhP9PN6E69AL4RK7SIA
XS3Jub5/kd+hzvPqRYyNcntPFjLm3VACElVOPfzTatd6XFKlksPxZStFl6AeCgX8
Dz6T5nLBJhPz8MCIiGAFgVLizRiOyJdQpoSqMdJV6kp56Po/2UYkmgLOEo2zAJ0a
sBvmRA7vWYt+ovH/qTKyabAJyY4UBNva8XSWqCrMCdtlwTPjOjuElaUrwrfbWrH2
D6sM0i7S+ZxD2RetDdddc4tddJu4ZvtMOnjYDW2U7GFolxr/qubI8iCsYFmeRv/U
gNYNv1raOQAUKh7SpYZIIAQ/oiKRYYME864y2n0TydTB1OVgLZfWkNYZFf24wtY/
W05+i9n/OsZUTOFayELwoCPU3IvfSkFfrXIJvd2WZEKEEmLWcJidGyLIyu8KbeRV
nmgjVE0wE8BAXtWRZNE+Rb9dgDoYhOI847EEf5dkaoQU3lPtD03EyEM8W3caSrv6
mnal28MPZLZ/LPH2fHr+lv0fU3KqXisoSYlDHvK2gQo+ZvwzYP9Q2P4mrrQjrvu6
qkUrTlD2xSqmWQIpt+jZWmJteqtthK23HYorhXMurSTUC3IcdeEQBGwgGOqZbYZs
EY1Xo/8sutK+IQmRA3NIa8oYWFiuxRT2qpn/NWqaNGw+rSrpfbEC4AF5l1c9XLCV
KkeGJnz4csIHC0ISLro/ML2c0DPENgYj00WgY9PpyeGK90zezG0mOthfgbrJqZtA
ZKASDJte4LZaJ5nJkhh7dae4as5R2j5efIzakNDw7jjp3EQfdLlVFinxAV8+HGwH
+x5rZJFLyFhgPQ2YErSM5FAbbS3uf1T8i9ffPaqEmI4aHV7PUqoHGBLWGV0+fxrb
iDF2VdHgThRiX6zyxSywhawaoraV3qN93R4fJLgMJxkL1jLhhbdrAlYi8Z6jm3LG
JmiG9vlT4kXaMMFCptxfOY5c0g9Tza7CxJuzj3x3Av8UJKnHx5GnYfZlwdYd65ks
akfz+T3LUvextJWhIYni4B6mmMlJu2W4ME9yRj9rU7C5Fa+NYyqNTgTxl2hdXL2o
bedvyL8I7UbYoP2BroPuPHkjmJmV/miACe9FsUZYn1eeaEmlH8BJal9BaXajObaq
gGnwRXgfuXnYOoDZYRYTURfqyeJPp//+UvPnH+cs44stc1BcmnVhhjARdopwvuDi
nuxkXcNl4NAVbcnshx4zH5oQJCUsEEShDk8wwmKvwb+ETbq2+ZTgbY5uNSZNLrgu
bcvv4HSQuHX0Aa7y24wdGJRvIXHxYclfqmmL8rvkcY60vLghn8jIkOYTo68c/GIi
T79wO+lUFu7uJ5lSYTSTV3/KbOL02iB3POrv6Awv1ZRsJ8QEpYkn0gi1J3FuIirc
Uan3h/OMw5vYMsnzh1vHEZW5jBO230wBVFveAVGDs/CLUEKYCy3l9Nl6Hjs42DEH
jjwjakRE5ev2IHJ/CuJXhJkmGlNuxSiyhM1NDpXORcu61zJRup0dnNwdgk2S2Bvd
3+K/jB/kNuea2hAJ8WwaStT4A/I6INl4msO0/vhVOfhgUWlhnBuzZhletC/LfvJG
gX3NKtjR2qsYxtKiD1HIOUwnszmFOQQ6NGn23In+eEBWaT+pMPAVYFXTSmAMDtxr
cIDzsLT1eld/X+kdI51U5iZiVDUs1AqyRQVGl3gT4p4wvpdL/ZzjSt+Gpv3LiR30
lvmZdQE3EoXLV5iZuTpYeVmfvdfW5y7u6C46r1JmLCnPngtgairVGYM7RrBIgDrN
EwDmyLzNkMWkDJeWsUZ/ZsSjmqkKq60s5TFBfX+X7Q5xFX6W4z94SKFrzcdBPqNe
fYl9Pl3Q7G/e2XNumOtNFDuOuLWKrKIk50P6nb9pv3I8hgToc/83Xr39XvM0VxsC
xqp7DCOyFb1bZ9WCr8mdC+cWSDsU5jG40GySJVqlljQzfiI36mjTYeHyA77pHYN0
albsFxx7QCsEUwFHm7+hoRUS2gR1cbm9edPqJtcEx8UUq6qVWY39fvIbWH3861b/
pnAryG/gC2I17POvmWnTXTLnOxmBK34dFqmU4sacGqCYhb9CAhgG1BbBnuWFeSJD
yN46zWd03fkn4b1PrCfCerL1Ai0rIBgfzrqKXdUsYESjXTFpK6VtUSJzIUh/hq7D
U0ElhErO5zQDGXOteCob8Z4GbODVESPs8hIbsJWnPXdIaxB+apJu65bdYiWC4j+R
X8wuZ/nbD0RNj+iFIz6fgp1lr6yh0lVY00c9AcH6dDXpfVy+Cw55aZKrXJeE3b4s
iYn6WWEG5L2YfoRzO/uE5/c4jpjgr2kq72VcbUf181Efjt0K8Rd8K9GA4Ne42Cm8
V6V0FTe5EdRODTaVAee5qUqZjw1MJd6TZcfoNJNoWGvWbwLrU/UZLEGs4RfFpJMv
bsvvJ0TwQ38802hjVFY+qb8BUE68I9CzVGPb2QNfW2ur3gFwL5TdgRUX9lQDJU7L
bL1wYvW5sgK4D01oQMDG81rYarhbWq0/clNV5gTrSrRH3xtEFLWfiEjToBCQ0ZpI
3b+GEC2eyt+n5Bv9cO2pOTfywwQzYYF5NRFEiW2WAWEIs8WLXmOWcQYYvl7fhP9a
UwI4s1IXKGVuYgO7EeuDf3z0aqP7xsaWTIl2WlVuB63ZpPeHXVyOKAoOxsc7XlCq
SJLVDfDQ4WU2Vb7GmRbpwnF0R0sLNuYVyc6b+xTxYq3JyASvTkprdYDSJoIdS9ec
VjUSUjeZHP3/jWyD3qET2moeGJt89JUNZrP8euFadQO8KEh3ZtzqNfD5dAaEb8Ae
Kr8zsk6pjKZr6HEZKNl2mIphptgkl3WXEPmkiS18hnuMIHE/iTVQkwbUFwERNxzS
AWTWWLxftjD+GicFWniBi8iZVbMhTxX07kkEteA0OPA50aZSaSrJj1XFCWrPxe68
bttxKMkzhzhQf7Z0cKvjEDSaiG2ZxSvIZaKxaAzkC9RqIpx+7WvIWVeeu2ASxH6j
S/5/KLUd7LjveYa5kH3UjdAU6NEIgtjsbhvZUMLZn12cH8ol4CnfxzqoHsyXixID
N8nB43pZaWg0W06GbtTyLNqzNJxdt5lGQuz7ZP4ODz2fXBDGN0egx29P16YTynEI
pBGAUdebFkUl9Y9f8m1vibsH5PHonsKUt4QYwJvijtZUPyQkOQZL1nH546rv4oU9
w0UxoHYNF1S6lbgk44wfWrtatGyynamup4mGmzIeAtkBvpSSKSVitH36tnE2fwCO
XQon47xqtjuRi/0hOWPoV9lBCIY4rsM/1TlPXqH7JUYmkwqHXiEA8mIUK2+RQo5V
/0zRIDJJC3QARAXc+OSyVfKAGzPimhKXKJG2zn8Jna/yfAXRAVYLyJLnZaf25su5
2TvGX++8PQKH7x350buCxL5if2DDZBcmZoGYA8G9QuInq5VMOYtPh0iNdvzxP6wR
PI+bbRxvsMWjjpAMELuhUfDGCV3+WFcTgoqwegz4OJu3kRBJACNqRLSZw51jmTQW
S1okiz5BQuv7gWgs7Qt8xNbeEr6P76QNtq62jJOAxgdRvwqve+8Ku3LVMHda6ALz
r+Z8NtFwGXgMVmjZNbW7rK183uKptfjnMBoaMMgvx3xTWv72yCF6sGUAJa6l6kH6
/rzvRtnDKVo/OdynLQE5+XeqxxYkGDkJv4BeQQ11r1PK0K/UMAPNjfRkU7fRxTmH
hePWRTYc1LXV/wCnGtbD47/8CLc0dgCpnLZ1B6UB3ZMrePJaShQD2gehJJ5iMEK+
Y/Z5F/xeUzrYNAPBkXkk2E8bWY4EyxONNyI3H/3tOLAP/RluLLGTNs8EW1WyeKXm
1jUX25Ltn202iOZcRtXI3tMeMBSMUkg1yPk1vN8xXIenaV2N3Q3AfBNshvnTGpFy
oR8h97NrKI7l3Dqbdu88Xol1izvFZCi8S//SwtsBV3EML+shR8aWs9BOgOQRqm3R
Zn9lrjiZkh6Zq4tO92PmtThzxXn+QcKyaycLFZ9hDJ7NLCT5Mn+aWDd7l34Tc0uw
g2jojNzYxEk5U+bIhCYdVFHLHmxraIRNqmOtH39gXzC9ZuPn6KYHpZYaff0Ra2lv
5ll2sjBObcbWvTE39E68qPiHo949QxFgNjgAlqf4q5/fD46lzD4xTzD1Nkffjzyp
Bab1ycReEDYDVKJtZlFsY1vZVHlUDVuyerIZia4QY0IUyR4OIkOQV9xgcVKoVxJ3
YeCcAUOTAFvh38CURXP0Y2aILVcmGAPreJ8l8Yigan3nbgCb+9MCNhdUihkRVvQE
Zo7YIEf50CKXgMevEm0R+Jbr/d9Vl09i51ZJLztkbiUANsJ6gBd9pTVSdQzgoybm
ws12aIPjxWhBFzEXOjYs4/hvB4f+tMV3Qa3ACXunex7trUdtCwj0256GHBN+e1Me
cWvxbFNylOl6EHJIWwqMQIV0NMIm9hfNZC49zXwVcqITraXrpIlsUrI6ohWLORmB
NsRZu0N69XfSkKJrqpqLtCkFW6MhwmUZOQwvqL3SkFtji1FMN43B739bYdVx92x8
Tn7T4sqVGEuqHqdtrgAu2sMlhQM1yEmUXoMqyO2KzSwe8l/e8/CHccqv8G7YO3Fa
OGDeYre2DGaog+v6w9+/fMG2n4lISMqG5q8UiHF6htnmHY0X/hCXengkTz3N+oAV
FsvkdAGwhsXqAwLrdXFYkk9qVWG7Ntkzq1QgilLarhDfCTk2vTffg4Yf1lxVZZff
dSflupRoJ0JHjDq/Hw5/tEBeA1Y3J90MjR/us3cPnewgwCjJEMoUPCrS1zaq/TYU
7X/GGqmTu4Q1kPFiNdP7XGi+aEazRxBW9WB4eXdysK4b8fQoDAitiBO7BxYJYClA
d+jairXc0Qj7au2Y1TpDUgB/czxLGjdBKwqBuGIYV9YcJfTVY9h74cF9Ua6NOxgI
Yt6s+jTFH4e4X02Ct24Zu6PUBEIpNd8GfLBnMVj4ev0r8ywEWKqXq8cmSAo08F7D
xhjnv+8BOeC4OOx/AfBdXU2YgccIEswNfXKHIz7D2tD+bBkgg0a3AkHnF+feiG18
qaWIbcRUNKG4BaqiLkhonbLcvMU8bRd0x3Mmnvzd1wURnjyxUTbYn3bwLoUWSiQq
PCzoeJRxcGzP4WNcY7z0WYM5Te1UKn1S6T4rITsMklD9Q9I9u5cezkg4jktmkNF9
9ygvNg7Gqh1Q8wstEzgud7AB663wMBNC6KJznmpAI2z1wp6mx/mh2lAm1lWI1RWu
kknU9KnpFNbB+kvZs185mcXoEJ98FkVKCuutxpIpHcsLcZsXrpXjBojP2+CeSLzt
iDk9+LcLa5zOT2dRxm4M80XrqzoKGqSIPHtuu43NiG0XXbcyjVueBGZzljIMh70F
8k05gIH3IkOhbBl5tj1PDQ8Spf9xxhAkUF96J2mb7j8LxiCNJenamAZk4FrU/sxw
qYGj0AYW26BT4Ao1enKKI2UdFImipZwwkWIX5oAIkp2RIGbJC3mCBaPszqeZLPTs
DL51twMYZ0k5UKtgJsirQvgDpYR3fAIw0P4sIxTkKTFrsZ7EaeZ0768oDHVVwhu5
1XqhPXUxUAaodEH9XTXgh+vbcw2wZgroQm8GMIVnSJt5MVI++Cc9chW3Enl4T8q1
m37S2bD3cT2wiH9jQu36ooZh/Ur5AjpbPquCM7pmlGIkPqBc5s+KNpyNcgmvWlpv
MNvgGVshLUBnfdAu/gK4wYNJhvaKPkFk5De+y+WDIgs89hIbj/ztTlskZt7palEE
fPwjB56jrCPN4CZI7j7JOWIMIL3OsKjtDeq/Ubc7LI+9i+OYRw5EwWL3S7sZ3zku
UwoJOdU8Qb051L3ihVturnPaa/6zcmb9VJGH8CGkIBA2b7P5/5R0djhWt3qZgTBI
s9VdPHXDg7UsVddT/JTUPftYkCuTzfvFPAudN2Yc1FZ2v5buRVmrzjVXikwHTz0/
cbArYFe0Tm3LaO31RPBqQ1ZcpucK6CT2cxLhCzmTLp5a5W7jDjvW9YSpA/bn+Xi2
jQAarBxMyFDL1ItdW/O/QDvWKI1j540JuF8oBHTwNGz0XHnl4uVLxLANK9OzLBmV
q+sKX1KL64Y7lSyfpSmogKmstawr92Hy+COxmwIrcfirblkAWRFbZo9cu8oucKim
4dSw81ezgYVMFWHN10WNrwpYgx9pgc3VDjGuQFb1H3Ri9vPfqqIRVkRCFAG3hOQi
6P77qGqh1+8dCBfx4ALVDPJATRYuj4nj38/0iKWSpB6i0gtpQXCmCTRNBwtDwAED
gXKsqTghWpyvC8KYwgEiNqk/b+fUhAyrhmsPu+YGhIQjpmNJCAFjxw8juUbdyp/3
7oyquvIBefrb5GhmFa8NeV1uN+t/X8KEW9YXDNh0tISr6DO4WDewmEmpD0eGy5On
JFcUaHWMIuLncIM5mchL+eobV72Ij1bztdYWGtsZW585YMdvkqAOEpX9p78Or/wa
FlzKa0zph2f+fXTrdv614bpJUxOGBEunJcweSDQHEoV3kiyzoqrcPRiQ7dFb67QC
TzwFc3R2KQkK7sMG9RuesHxRMsxJlEckTqaD5e9mzYbyEpx8Up2t/a8iDyuF5Bbp
J7wPQxu+5DWKq+1IeHgmh0WlCr71IKxXi/X0HjSA4Z13mxVbzk0t78Ytdij8BZ/W
SeRyR4Y3b6Dw4T5e7/4kisjlrTfMzA/u3J7YGIJTurhstwsM+mcmTYPgBdYa5KZT
BXVKh+/3iKh2c1hl8adEraqbShUWLyP2E4piZNxPXUroEEe9nICjHHXJtZ0c6lSX
mxSNzE9bYimevZfWKnhqNXgDLU+aUPOyQZ5s65VIp3p131L31Av/UBb4/Vpsc1zF
A8D1PNBu50VMUXdcogpO3UpJKW/CzVMlvNl1o8I4aBUCYdbd7atZgmM8C4W3p2Zs
6i5B/7zfc/e7LQ8LKrkABvGd3tBKtXvWCU2MnlH6kfNZ2NXx8cfw+I/m3gOT6j9K
BKFDInFhH2atvV26wKs9NuT8HDH/ZAv/E2d/+4B9c8uPjndCbi7fr6k3vaSqekYL
ZJtRPkQB2SadqN8wcadjmcNcsK5aHOn8lrNyFOcqHJ8M9oqBuSvipCGDN9QXrP3F
3Wab70J6BCs2gcUIRcI0C+TIblZehiEi/BMuO+jWqciwrpWbf8gLo6xc6spa2qfb
D9hT9Af1DIQLQRvZS987ymVD51Z/g5OOl3iETK2YKATo0MHcT0KqAgIIqJt0+mEf
s4FrUOnW5JaLZ7oFbMZTyLAx2uijcGR+noB+2WX8H2wSVRkYGfjN5bApTJ6Q7OL1
vv2m2c/uHnBu9rTLTV76VwhuPCMEIOk2EYYjQT2y+Og/Ey3DY0FbwMWOYpZoKr9b
24FNAcY9sxBzceXqDz2ZG+nYOaMA5ONwo2kcuBB4dfUZZa0ebpkpjj5WzCE07uTS
RSNdc8Cr9En3AsZ83ZeUlTu6ZP0aRPXhxU7rR30McQ871RnqzHpnXeHzC6gGukbN
rA56mtGb+QSgNO5gTnDtlwavA6wXvYfT2vtEe0u813nr0FAmAhSrYjQztkmMxQnm
m2DPPP6XLg4tz1K/3O/nruvhO0EINOez/+Qn+6lctKPZW+mG9YRoKcTgM1T81DCG
q3T7MyGVP+ehi4P9gbM+2xTh5X01pZb4ekZXPoZcIyLRNv6wayxvvFxogoA4BX7R
Maj9BQ3pXNmZm54uEIIkfjUCJsh4HiGxqPdg9CQjvp7nf5i99vEDIaAfRwGhFsYJ
IiuiAfvMoXIvDoB+svvmE2D/kTP35o5IAOK5e938+fK497UqwFiWHbSX0j3J90UL
ObS25EW2K1fd6Ohg0y8YEW6GyfxuYtIOgaObGiEHIEo5RLk/6VGgN2qo54S2w86f
m6kkfqSJn9OxnDHjaUx6YyOLtViX9LFbAuYLkb7htRtSBWy2vizShtJ3rJcO8Pgn
8+XaIdFKQ6TGrd4YoiPkbBw20wMeKXfDX0KfOSwJjJgq3ToLSzQhjg6jcWeB/47U
uZOHGcexrcu/VVfrqz2x+L5JFaGj0eDhrbHdbrlQfLQVG70cxoo/N3CqOUMOcz01
8Tzbif6+k6tOp2gcKCNyKQser+tnmIsV/+D85y3KzwOBYh5msLS+2zU0cTsC6lff
TRmMfoaaE/kbxI7keZNcYhFOxxU8oWEpf448rzknDlTHki9Y3NY/2b1vEZW/SIhj
haOaDL+MslFyH/Jhai9CoHCKW02sTU7j6z3hBJ9Io2eomH5SAlnneNGDCD1Gs3ya
HQ4AkS+pps1E6B8rlnPuZFJprz7hUXNG3x+nSvK5GllWKUh8G7N/hKh5+Y6U7FD5
sfBRLpFFgRmJ860pMUaVE+lbnI471h5xMtPx2PgIY+7p1lhnu0ywG061QENlHMSK
hd9bzUgxCzpWr/SVB22XzPn3GL/89rbl9CQ1C608CKwzXjLTjREwGN3lu4S3BDc2
LYJHIouqw+3unegW4FYHuJrGGp8AIaTpgvC1g5bLCxNQ0r7Edl/hoFSRP3AGu9Za
wXLAOvIIUNaJYuasiYfUy97ZfWLaNpg6WevDfSiinVjLt1gO5y0HVWQykDqfVOhz
L/1aZlqNOXGvJ8iGk9niqqKSzd7P2bICkKr3cVja1Tk2cYE1jcNN9Li18ddqxFhS
zOGYkphlXceVYJqvQEqqvvZJh4TUsS7UbWIAG/M26KI5eJKlYPdE3M7Qf/Fz0Z6Q
+GdutDktAum1xHRBGIjOosXt0u17LiGzwhBJrN623LBw5lTRxVAxCalUx1QtyYUh
Hjd+kIL7AA2NYM6GNpE5ctGAWuuYhtPkshjrXZig5yakQ+hzLNrlKb7cBKINf80u
Wy3HlV8AbOnuZg060oShqukMKL+v9GaSENh8rDjEWfsY4MPmX4IqP3J23QSqwiyO
rjYmZ9RkYsICqkbVDJI5Q/VVuCLmAJ31Aup1ogkG/eux2jMylLMICOCm7tvFzdwe
KX0QwSKR4kaYJcVbt5wbc7P4XWKX5+AfzFd669rb2pC9lQqA5YqOtxWKe9Q1jw+O
P+0mmYjCNCBMTbdROgyQLqLFqc8YJGXBb5EddlS0GW38YChKKv5yhBkYNkftKrZn
s2aj8Riws5OOjX8LoSI/S6jq1SSrxVZcuoFDZi2BocYuCMyzSbFI6isXrs2nzZej
Isd2Q7nWh87o1PfmJsd7mSfOE6PLdPj7wz2ipLiQ43S/ET8sJqshxlZohT4K0Uh1
ydbi6mkkNYjZDR0JbAmWkymOy3zLmYqwkJpzH/PagBNr3pWD4JbAck6wtOWgPL35
876/Z63okrt8osbPj+PwGpLD09CxBJ5lWaHG9704FHNBPin9fI/pji8fUETHxg+M
EL+ASOEws81UiNfVnlHKoA02Zsmv8FIU5SCCy1LLKBKGaUoUlwOHSOOpgsCubz2O
JzfkAat92qKQY6qRGi9dkndZbvDcT3u9Yy5f+o3AcfdR9Ayv3Hs3B1qQaeWS8EhZ
l+PsWAEAZdBH+8iC4WJ+GfQ9qssPVCTfpaYuAKQmAJWvHafiPX/4Hu4s21b7SBoE
hJX1NSOLDmilyR+ZJvlLz5Uj+Ndu7nYpBWO9gP1Xt7I5XwEstqLxCtZEDI5oOC7q
lrP595RoTVQiYlotf9O6zboG+AKLgc9Sob1izkKAC5uZMWpovKC/jUwidahN5n3H
VMP9chgMKcRNM4CFJfTWn+MftGY+llbPSkxHMFzFqVaJ1iy6luWVWBQoVhbEbJv+
MadE3oH3vNh1ivRIRdYZfBmVUYHectTUKBO/qX+MJoIzMLhqxfmaxRn5MQoQPRpJ
Aqq7T6A9X2cMdIrWU3kcbNp46oXfKx0a4pC+GE67QucZ6t6/WObAIPymnCCHLNaZ
TYcRk2JFeiUJN1OSsraiaznsvRK3M/OrFznyIaYm+HoDYADs4xqk9bI87xk+vJO0
4/PCwbt3fjUDFInkgTYLjiHikqvnQKkWVxgtlGoDFr5vOTti08vs+ipizRHqpzHk
FGek9cOL7aYxDr6X9WqjxKg43LwLqOrUi6eaEPNcP6k9s3/XCiKLblt6UZmJnqwD
Hr5P+gMYUDSNlDatYFsGwsG+ALdbnJVWKblf+0fthPxa1hvK/GC1u/tCenUqAabJ
wqKAkUFMwQNgiYui+r68UrwnIHMUsKcJxmImvsdiMx/fNnDrqKnG0GZniy18zCEc
geoWVY7WR6n5ZMoxUCf9HEhS3MfwfM4J5Cep8byjHha71V3CCJuphxLaP8ZFGQkK
iUmQO/xKyUOmlXY4hk0pso08u2Wxu7Med5xHlRv2TYRbnM7fsoG6+OsaslzMW4cW
T8jrLOatIQs6RKU15iOB4ieLb302B4MNPSIj4MQwLAXnF0CW7OhUzOqlxikMNy8W
y4jsJ5xV4k0soosS3EIZ3hWoDvPxRUfoItYU9AZPhHqvuTO9d9ljIE1LPd3cYvJb
G+s1XE8clzaiIm3XmI8AiJMeB3P1Ex1yF284CB+Q9aSgHQ4911v9s1CVmr8tOfEE
RZWVYrzLRGcYwT76EFoYDTTw8WhNqt7XvUdUA/OOdZdH705DcQTit8j3RnNijwRR
Sa8n2z+zxtJvUBhQ+/dAsJMIE67r3NTfK3eG/Ojw0x1PTEBmEPkz35unpnQp5uHn
SqQudV03ZPBNJHU2FQZaRSSP/ubBgHrM8qN1QW9VYheeDt+95oFR2yJdNP8GHwiI
be5e2HGJ20LLEnIZSXVUdbl1n98D5dLr3b/ws2VISxMZkGrwCVP1RdzOiSPFqP9R
uJgLlZpCU1XF08N3u7r45AAmMnHDsmUrfkFUQ3v/rLknRoj/DgGNYe7SrDPzRnJ7
Zfi72qLuQV+65AJFM6Dm9Pga38TMlMfk2MKiaRcr+chBylMPGQuMSc45F03VSJbY
lkbr/2kb0YNZkcILGzi41xUjGWQ+u1Fo75GdtViRsFrAg9qA+1z5eO5EqbgSYszu
BdP5pb9T7Z65BcDaQqDL25svkc21yjtXhtRPMN6RRh08szrlC9/jTNjBEv4jukNt
N5mjnWJjvi7fLqNsI1swC7RSe7IiiqYQyfXweuicCsWr8fIKbaycwhiobvEEOnKG
BVLczCH6c0v6hqQyFQ+urNPfAplQTlMy0EcTWnR+3JQkSvXzTl6HNv/TICQYSNK3
iLNz1S9DjlJn/LvPXUBVvJYUVTFOTeJD4T0q2XYaJQIsxP2oAF1Bp6hn/TPgioZc
pgVhtWaJZEMjwRzQL4njyAI16aTR3Hr1DELc8IbABU/L3GbMOTCiiPiB9KlXexx+
kzQzU/MuIelXWpsqOr892ZSJkPIpXIv5rzI5l+xi3QRRd1tQK8+U8iqA4jKtXu9y
Kg1lhdPx3l8tqDBx66LzRsnjLwTF6aoaKeIk8asPQeOKCrpK8A7lKeorkC+H9QP4
79N2Lsg6QOR/XURDcYaM2bvjkARq39hhZc+pG1vrrs848E/RmKNcXrxyX7cTvYFg
PLDEjEcjPIlpM+UALz1Zf95xGqRKGZuj9ehbKQSAo248GbjnP+xHq3OTVjwvSGRo
MKpzRsBjoILGtq9QWC1zp/7mmSkASDUPZ1cnW1/BGF77kVDC9RyY0K5Lh7aMySum
ZxCiPjX29Xww65awNK/cH6C+UzwM52sZKuCCh0k706ZVlwMqfn4Hh5NPBZ+XIiCm
ocO/vYeO3fHzVuSJxpnwJgjCscjMAF1EfPOfyDRHwFstRHB17R2haJWy+ppuMO7K
ygzmt6zc97QrVDMeK5BEDCCczwKAoquE8bAQkyXdt6rxcDV1p+zqKbRA+3An5LTs
VPncoGOiUuuiFpMzB4vZAJysncln3qZ8fXhPYmDJ+lVPQ8F2OSqIvej11bXj7coq
8FRjiAM8gGw/5TnjPbB1G+7S853qHlWJXhiL+Q0HhvB58Z/Oc8rtpO8PpwyGaqEx
HWzhhLqg/uvhSo2Suf0R3UXupa7yCnQyiarzp26HmNc66Khwdt2GhEnd7uwEDTmW
zMiEbJWKNMvCFsr7f+rfm6aS6B39SEPTVtDrzzLb711leHQqXTyU0jmKrQJM7S76
jfzi9rFvzr4rfL6vBkmQp3sp90RlyVRkArEAUOmyq4JOFrRzmtQxdx3npWbSMF1g
eRy/vsiwXtsROZvsW3y2IsU7i1zcvRPqMbhUow4GiJJKC1Mjv/53OW7PjgltNxLH
IzfOIbj8+WzBgVHVveKjRtIUi/X2MJhJYlERYReMK05lx4+NcpPeiEvHtDjI3i6V
Dj6j/H2skwdSpCsQhAj+Tbdc9T0SD07LZSV1YDg+SgDG7Tv5van4e9Ap6gEGZ34E
FKXRbQMobKITSv4Q/kAemlVETPRlCU3PgQj0dJz1/5dIfzFCrCVmo34EC3Pwr3PB
tuQ7Dom8kcR8Qn/2iIZhDIixsFKspHvL2bz2Uiqmvio4WxCVRjcyDSNgWlQ4gO3z
Wtf2z31zK3thE+tTya41J+0dn09POAAqL3kPqTFVXxWQJAetMnL99b4n7fPea787
dr3pqjJ+inm0BKSQ4k3QGXP8gIULkk5zhB3JLXwDQzJ+BNLwzHnAGAj33FfoD6kR
eM4AQj/G2Aut1Ait5LChsxe3CAe7MTWx2rmYsC6eUZznFkPPP9T3+NNs73WyscOO
hAtHcpS2AvxDn5lq/2XE2SCu6oHt8nZjr2ifQNVEgBulO3ftccDpetxMMO6JVKKz
fl+mVHIkYFcuETz9ZRRCtTi/mFlm3v34jToSR5yVNvwiJohAsfyZ/FvVAWWiDfJ8
KIoLhK+nrm6ewpeGQ5uSdkWtLtOPl2t+RsnCsTxRs4AGqkRRcjy1/8YeZYYOWG/v
37XJW/8b7VUrK5ic4k7Q7gMlCAfstedq8gJ/3nYum8F7vuDy1EB9cDd+rh6acRYv
lRZeC/fmNsNKkVBcMslYE3TrIg8Jx+DrCrgiQ0r0WA+4nsfAAbxN+lNSmvvSjZFM
iQAzNBdY2QZ8hnYG29vHEQu9ng64AUBUru6ObnoJUxiFX6e5CnzEsfN1rEPaZvLK
ydpKJVK85qVhnhJgv2vw6ZGGo3jMM7vxyNrKipDSYOhql/BmqU4yPzHvqFIzDKSq
zBj3GVSUYGxtbIDWzEHpmAuPms6GQ2bOvEyU0SYl0cpZo97qWQmeE9/CwJ05Qut9
N5ihab9yTc4JV3v3g+/R5CkD2sWs+xoeEluq68/ltwWRvXR2JrNKPIHkfi/0mcsk
4dP9Us4xR/EcFbje35eLOnidPHc4mlI6GHdxTqfcavHRZrQkUINWewUCxintFoUu
3JeAIvmqqBQYb74NqiTIYNq/daSkyn+z8lNmrMVHg4EyTCioPCaqVlK0e3/cEbRi
87FzHPnhTOHYW3ADsmacXcNIZRQfaM+9xE38V86T0zuYziElyhvlCwUFvNNt7S76
2nmC7M6a0Ctx8JvQcgOsNEzTHrZsaFQCvtuPZ/wJoRcJdHBiiRdJU8RYghA4CbUK
OWArm2vPdh+JJflZItRIbrtO6epEqnF5PM6r0WT5zHEK+9iSDQ6o2Kqg27xcBYvL
yE2OE5grka+ghB9kI/rktOl6RdR+sjC7/IyIJu1FRxoosGPWuZ+Op0DkdBPyyBZp
xZbiKoEaKFUnctyWD455Ed4FHsTbxWaOsj7y6V9qu2HRCEk5pWEpI67go2c4fmKZ
Jsz3nmfJqyFdx6anm2eOBVISdqLycTpDHaSr3TbHPlGPxaBhBDTCm0sDGxeCvM+D
bkP8EnUHv9kmBdyt1feaZPqetjGrd3AIH9nhrckxI0OBkFb22dz1YDjzoqaYacPY
nN9wN8ZNWFIICBOY7iyOYkOihCb6Dv9KyzDcNvyPK4n4cyYryUIkJ6zqe037IzQA
DdwIKB6YYGjZ1yUG6PM96Flh3xqrVdRtxODng7EuYxkLrgSHWsvA5jJa7tdoNNUa
Qk7NTfg5QYKIwMnQ9FzYZychz86mWhJL9a84FL+VJiejavTFMoTsLv1gW/5esQwC
x4dVwADAMSrmQuPqXSYinQdsbePVWLZgVAKxFlUkSuyDslY2TTqWl4jG+P6hXiJ5
8JrL74cJRJ0v2AMFVhCds/WKST6x6q4uufequJeFk/JKKbnDqqYB4N8s+Z1dH15G
bodZluM+JlRkMuA1lZsOanJ8POROFVLmQOZ4/vofyBRA8erP3IHSDtAVdClpoehi
OVpF8tFts+wtMG5qLbNRtByc9OUtfo+DNNdA5SyAhYJ5zpB1zAamHDIsRMXMbORW
2tfrtUXSBLUgdAiKEB08he4YCSMNGsr0381IIcn4acQp5P89OZ3zb1atdLTwP8yP
f1rnlK2e8ub6V0Fmknt+vXRtNtOVIVKH/acGiSf3HAVadn137aYKdl86wW2sFmIv
N8Zpeq6XhDwtR0KDHf1D88ZIY0mbnWjlKM8E84UDJB6AA+eHK33Q68oeOzdsaNVR
mehgkfryf7gqQR4EbaQk/KtJmucUBZLdzCJDmzJu0CjX8Ci4uNvOenTmmjFqmVvu
sEzD6T2E7XuXusbf/oxU7tlvaOUUH97pSDQG9rFBKlcJpEUq5YdGk2gAhan9xRpa
ATSdrr8k9KMvQTHX8+DTXW1VsAe+EUsDooW4yfNGs7j4WJ24y1OCzFO7iKP0GvkQ
sz/GqzgnqDwjXU0j63u4Nx+2VZ2UkX7nazDAvC8GTtwAm2qLKnjeFGKBUwfIGcG2
0nrLN8M/5oCVK9FWs4jFTCjcvB1QPiMGGluKhnHDB9rFqv0nv1tE7tXl/0YZ8Ywf
ZbhP5ytXaCI5p9JuzWpoTYdsi5+1YEN3HbnNczqIhKDF9T33k3bVV/L/K5cl16aK
AjwNrFXGFHuyVK2SStNCV/hLEO2C7qo7LTBH1telurJWrgYjlRH6ei7VLK7CW8nf
UG+OG1775w4QchYr+LnJzrSLUm7eGH+oiwtX6VJceJmg0EXCzfINbs5dI/Tkp7Cv
Uyq9JNuZsRdj5vk9qwMKRVgD0df3hCpGLCrPdRFKwK5ookqoMk4wWnNUh2vZBO+b
wbH1CXx52+xhkJ+e1g3AgtW5WUO3UkBr2JuUIM5VRK6fat4StejmbBMduuU0X3I4
Z0XTjd2M6zAU/CZKnrWYChQjYFKFlMiTZ7lT1Nozl9GUeehRafvBuOfzRSu9P0bO
PD7N761AQ/W9Pwqb33YzbLvznrRe2ZaO5O3P5in8Ez7yNKR/zbPLQIs3/VI28QQg
6ZDs4EISykc/kAPT5AqfVUFSVQcrvvzIUC1ZwMxBvx/RciinJvUXtr7g70UJetg+
Bh9ZFEsEh5ssn4okujXVThgVtZEaYk3cQuJe/ekDUQkgZrsq4/iU2n/dnN72ro82
e37sqlkj6HZD7W1u0G+KjxEbS7q6A/pZeaU3uTVRPs4rn9my67LHdeNt+vG29LAO
WnV+5xFKNfdrYPIP8pcUXWMVySSI7lWj+E9X8hsnjW765UhnVo82/GdMYNrTLDxZ
4tOm3VljQ9rDFm8++5rLktd8b1I8Wz9fIlmai+ww1Rr/5SUXFbeCGywaTvbJzt1o
+2Iz3AFVaVf4DF5KrmVbhrPS89zxXov+hCL6Zo3btthuqdHFPf/siPQzPxYxxjpS
rPaCH1YaetbKrocU6pG+4TqNfSYqi7U+f0/r2wj99zpJenQfp/an6gZ5ejLkV6y1
euUEdWZ5aQz180uOYKVPYIESyaHAmYpu3ul2/bHQK5clkZvQuOcLB3iyQ37ls0Zx
QsIwbWGNOr7TsGc9kSwd8CQF0Q9dYMwl+udRtYepW7pMWKAgPux79K13fCVWs0eg
cVy5+zgbO1ok0lCzM6MIKSIiV6vJH2Sd/b9Kk/5fffHkbTtBUmwfxkAxawDqqfKD
qeRa88sC84sEUiNGqCRLcZ7vzk8AY09GCpsJROAk24socnB1VhUi0vc4m8oC4EHO
hndomln3gaYsqHNgluU5L1DXnjnhZNqb49imdhH/391AocfugD61kE4mtxnWNc71
/MHZjUO2SCVcie+UYq/D4norHa0O3xhI+A1ZtDunCCiEg2t9YesiiwFZzguoZUNE
yzbFJCRT/37EjvLTYoCuKMtZYOGTt+AOgtRj8qiaeGvB1qEptUKTIN54FaRUzdAx
b8h/TR0voFFZAyK0k31z+Y1et2CCKqZVI6v3ZEHdjQ1Gf+WiG4UIYZD8JjuDAN5u
TcAwvifDoRZjgrmvXGXxty+/s9VawE4PLsDGbznjMqaJFLYPKIbQDODGZceGqc3T
3+HJO4M0m0ik6NurrDZB6Rzpikfhwi9Q+UcqiQSA7gApySHYfbuzxZE2+A4NDhkQ
fw/rUaHGLJ8JWs8lfen8xF9V0pmJAYHyuKpNeE60BcznLMVKUWrbw4DPyNijMB5Z
SBxh3MvYHCfE0aEXICgii9XHWF6Il5ct1iZOp9zmjzIKt2QYc8OLbt0fipISbO62
hGKqpvG292rcgEViO/0Az7noP8GzoPwJdHM+tjWrtO6ncgnuxcViXS2NJ3EhS+gS
nvPCDqUcpjAGQe2UvsXVSRY9euY4TolMXn06vhI43/1acU84qi+mkxJsvyKUwDyV
BMnzMC3jaGczAD1Fj2uUM9NeXRJY/wJEeM7nLDWQ5cgeLQ8/eD8+mlKmR2SGD1cF
mtHC8MNJhrCAirmfAGQ3hkW1OCzORA+qxL9N5GvgjLuoSdusZGb+XsaqzHv1uOup
3vbcLM7bjZJhS5WVxP1BCb+ShqihWkQLhA4bWJeI1CVLFAU3Vr3DgI/3qkjGzpMN
yNQ4idLOnL0aITxxPwqWoH3rdyGGVC3ZsZQ6+S/DBVD6TlD8sQc/+ZffSu7u7m+y
Ld2VveLLG9qLymGa7DT1Vm0HOgPN5aMEK2PBf/GSgHh3aWFDV4EXRt/ZilwIiQOX
StnE0WAqVu8yqbMnz/FQ0YTgOLBBc8XiT9O9RXzhUppsXHEHksletDVx4fOD24f1
QwdUC8emSTj1BfwCFrIwo+Gt0FVGA6n4mW/H2YEytYNGV3trwvz88H1PfJQmtVM6
l6YincrPZTFH+h9oiVQjaQrkxZvGKgmph82Rg/QAKUOQJS9wQ2h7guWIZBOctdmT
D04kiCdPAn2ds4Q8BE5xwFhaFHvz2KeQmMiAfbyC+VTzts/C4G6Zv+ATtuPLX5Lv
kPMf7b9zNkyiIU/Oh8kuR5AjMd4AZ5e6a411haUuGS/Les5MtFSJOy5UBoeKFIu8
gbsEmKxyqHDNcSBjwEHXcBDdKfVNgD7mg24J4nwObr1gmEic9oJA2wOxiY9VT06u
Xtk1rmcD3d8mAC+Hx464gOogmjwX3XJWDgpaS60BpHq1F+cf8pSKpP5LqtSHOBHM
1cXitJknaLcncmp0ngr1QkUm/qC1v9B11xRb4qD7onXcXzh0vQnL1K/sNjn94Yr1
NaJfcM8sxPbAxUr3oXC9VILYsYj59+dkz2EY12WBop5SfeCFX/rxlU9lrf3mrYfS
1g2tbsItFmkOGbgUl0TZ08cXReKayFFBnGn+SC9ir7gFnHHFiwAYDzN5L1+3Ej/5
4kdJlndYB6hDLIip4l/LCw+DIP0aknlO99APo77SKsE3y9Q1vnTD7Xw+vddIZH+m
xSciprq/necJU/X04eP1B9uoDuGWPZp3DZk6t2PfFLaEOg7E3SZySsBG/YmRQ2a5
Yrg4mfCnXT24S7Elvvl9gfhbTUmmUqxQx/wLpO68mUVM3C9xHArkQ9jV5DVQLoZN
JD9OSsxrebixNjmXZxX9AS1OubGqmGS6qdCXSNs/W+V2T2vcxU/MtvNBzMbYHffE
SeKB8vQJZCvBr/u6WvYtD2e2pEUjPkMGr6O+nQQcj781xjh8XXkg8OTP8nZyXy/9
14nv/el1jTwCVi9M9lIWrh/Ty9XG1MSYlBz8kSb3l2TZBmOb91q8rAI8vhJdOuni
akkYm/XSbetLEZRGS8rzihChaIgxnRRXYD0rSo2Jn6rhiffAS07NISKQBi3MR02H
0agfxXTVkUNxYmnJUWz1jroUG/8GnfXmKAQYy4xe92uLELpxPpkOeF0bm+iy27iQ
2sfpgTTKcj1kP/6YguEnWUzxDoj6jy/arhKwR4arx0uCVjIM2w1zdQrOxFsi7J17
Y9gr2+ssVxqRNnVyNqWOXmaW6bHjgNGD4o2OqeLU3vjngYrXLs2dAyJMttNSR4uE
VqjINVQKqJYF3Xtpy+bTP6upBB5gLR9qW2RFg4Ke5Oguy5Q9YD9dtqAuKLTPEHal
JfnaQOnHc8WWmQYA9cu/6LDLngHf6pJz50gtAShV3axrOkf1BOGc9ZvzL3c+7lLE
s2RKNAJaptxOY6m2BX85n9usesW7gGiOkzFZs7b7m6VOOSAtzUA68bQ7lKGZK8OM
+BIe6mARXuH933iVD9RqV/H957Q3TC1FtY0B2i5B5kBMFIf3WyrYSJy8Qf5X0dtg
fmTTNWn/i9Pc62KE+sTwoKQM4yhy7pDW/+mOnU8HQNYmiOzl3WLHnELjsicx1wUC
+Y9aW8WT665lSXvEnPY5SMcjCJbMKxvB2BJZo7mG8uVymuGWJTnChTgTZ50xrfLd
mK80OgDmslvfp1BxPKugdsuG77Ky65jUY+nB9gAl+Y7L7bZkgz7np8/3e6FRIE+L
Q8Gs0TsI+njflhs6BaOf2bx0hAkJgtgi/8zDporwUiqpG64uc+iotpCn3wUQq0G1
UW15x4GSMhcz/qGof1XWg9eRTPJwEYD0sMs+LCyx6P8oz8vD+SFiVOMLZQG2/ELL
yFazNzwWI1kRdctVuoOqjCY4vL26XarlSbFUGLcWnTPD4COlu+l8mLu2SOgumZ3T
flvQHldeHV3uw4CpnQH/DS0NCY3qrAPotXePfubQFzLTJL42zFwxVaTpX3mLkYHi
uVl4ZCrpBrwbLQ7vsDfDKhRC/W9S6qZ3uTJbZtuoIvnPIGvCOLXfnzJEI+UnlkiQ
dPKtM+atzFgxLvaXPvzoTjPDpkI0kTCmxDU5bDki/Vq5Dq+1rKarLLaZkP1Nlr08
mwR0slf7pyohunl+hKRXaIRk7o4ZR2gScEQtKkMEJsRIf1zwGdhz366KNYNVR+Wr
4PgDZo8PNfK1dnpDCzCqpv3A0i7eo9rv4c1kdUYL1hsJe2n/I15h+OSKBVQ+rsMC
h4JBV5tU2ALhJeyCky3Zvfl6UVwC6V17/VWS3NeFeG/6T9SW6v8wRYIAq2mMtbcJ
k0yDg/ZvB62G6YlE79e6nKOgiMmnpawFmHmtT848sLqWthq8+Nm2VlWwGOuw42WT
yNSK4ed+5XYskytK3zgqNjyGKbt6oTZV8eokEo8e/dY/p1RtUTKO1vYlH0kam733
iXlwQyPcvpPmFH1S85NYtTjPmHZ+JZraeN3VX8L8PJJrDepy88JuvBVwN/iBOq87
6SXXiACTwzfWyzi6CZ2nQgX/nsJ+8CRmU+1oM/KUGJLu3CVLOFWV7bNbV0UYfeHg
ZJMK2vEQv1QZpRC5EWIxLy7Vun3BhuyVS54aZXn9htaMWFZ/T5qV3X5sQIV8sIh0
dhC2iD1RMIY0gUh4EjAUXwT0oWRfSexylh9JJjIg5c6qbIQ6T3U35a395lCOy4QT
2WWtvJ24begauVn4TlxswqSySbB8oVar4e29n6kVagHDXmr5XVPRN/W+oABYrHl1
xvWwjHTej8haKuKKWgac4WyBFDgjG9eiAx0aoom0jECQmUIycijj+ur3OkQFuDcp
5o7JnAOZyONQQOudVaO/vI9Pu0bXkounupe5clxNCWveeuNQpXVfDWnrlAnETGow
MSl+zCFrvvE8rIx8mUsdH6xKudjK8Tq/sLQwlO8PrZkbhHRwjufKoQvhjZoj+m2H
AwtvPqe2aRpexyaAJ8zwqSNgtM5gryMzk3aHSeSB87eh/W7GRYzKaOcPFymVVwQz
qeDSmhHt6IKDtbMXNAf+DYHNyoKoafYGcGQrWODn7OG2ckR/a/YjirF2Tc3sr+jd
SlAGSOhTztEM/bxytXFbnZQnsh7CU+fARC5rqbbtLq7RO4lccnRwfT1CpYH5vPdd
SUzZre1PQruVX0jAG/AH2CWIo68L4WBksVqZq+7agvnitZuRPHpfilOFaMVZp7ZC
j91yfoFnzT72K6QLqAW7oWCDxjCfkuuH04vDpBk1OLm5TQBEBeJSGIX0xB8bpreb
DtYYs7Gk7ge6S4j2HmVXHgR3QF1GM3rlTKuuo0YVwbSYW2fvc/vCx8i2Nfs+wBEt
lVS2glrti7fwxVF3A8n8i47rPjVCDHCkqrkAoMXn0IqhqNMZjkoirc5n4KxAnu+R
4+uQoRgOvtS4O5u6orMOqWxxsqmHMBxZ2HvQE11Kq7rME5nVFCg24adIxHc5sjhl
XHkCZVZQn3BAW0D9OotgPd3VEdvReIEr2p2A9+dfGEURF7vXfmrQuqcEaxL42vkx
poQWl8J9Sn5GNd2kV8M11Jr/1RHSuQTgFEy2pQl3v684+TiMmbuGOulgxyxe/w+Z
0rU90OXqrMiqDySytU6DstQdblZ+jHtwNPaKzNSXaXmKW+D9Q0YJjKfVvlXSAUsJ
5t5sgou1XEfCEvPFgyff3X1qNqZ+09PWlNjHOVXp/xYEjyq13E+uhQ2zuQTS+bRu
Ql3tvchnb8cPJclG4CVtt9Khj65g94huSh1hRAdH6dadpzWySGwRGc/AbU4G7lqL
2fbYhHv6rSY4LNkMVuonzBdNbkJDLLh6yj0T2hF/Zklq4yorcyWmqo4PU8XekIjo
TsGCRynhztItKgOCj1M+EVsM/kR6eR0iurLiq6w6airFZmwlZ1yugiuXXdpESYdj
EW089pzEAE2cLzw+rAzC7ZmQJ0aCSHEdKB6rThz7bp6w3DMAsYIHERDLuowJPCht
t/TZNncNeRFhSFcLrSGR/Gki2psFLkVs13s3tsnZu8WnrR3MRRjSgU7d85M3FO0I
zbj3yvrjiF2toCxDcJm3UP3rDPilk+RB7iqo9jhK5dak/NrYnFzFqm4mPkVb6xOO
ZEjU+uCN+3uY0+1BVR4yR6c25CD5p9zxmePGNR1RbqErr7fDo0+Zct/DWfy/sZ10
M5jBGFhP3ai5D/inUPzn1l850zbfTu9AntypmLVNoEDLsnFrcATfj5Fi871JfUmY
dSszO7ixn0HKiQe//bl6+5ijDV6AxN+oxUoC4/BmSfU+v5xq8d1H8cmMfd09U+1L
9xTi8Hetmmc+BCqTfKBwDtEjX3dJh+Rl7oPh2TEGHnKejw3Hs8RXcaORF+AzK6+n
H3KX1TCAm2uz6u/Ai2KmWdLlnnNuI3igYdXIrqRPQMyWadmO3aNOdczFJbC7ismO
AY01Var+9cwVd1LPXJaRRIjZxEGsJnJJLnh5+bbDelvJPX+/9ytgVvq9rYqMdvE1
3M7/O8w1RbkCO4wbCiV3GXRMScnI+MzCaPAHZ8DumMcJmNvV7ifZwzxg8cswKgkb
lxMtHhhfa6UH5Pr3ViTdR6ZpZGG4U91mrkWZCnpT8q1xuIYHdUo3WU2L862UXuB3
SxiSl5P79m20HWgfmHmQT3hR8tNO2qRrKLCyRkh5O3bOBLyV2ydtg+RSKG21wkWD
uxJJ5rKWzzXyb4qtFNqMDozkfFmnbjQoHqImYiDM75984LKb0G3yJG0EKxDwR2CD
DpVvtkk51N7Jx9NBpRfEV8x/nsuKRTyJaJTbD99QerKiHdHZuHoCi5XeRxG3GbPp
EJuG4qeAypDnkyM0/+KjS9DaGGHsx38xTwc7Fj3kpuvLrjpiIb+MJEEDb09ZGYF0
kfBt9n076yBNlfd9cPJes6rQRI4zRfjuNUhvsqFgIgeJMyXUh0LjNJfjwBNlTqBk
1gDHg+APmU4Y6YTe//2hQlXymNbqrCuJi4mJuN0FyFMW5sUBcHwp2inS0942H0Eo
tNTz/kz5HmbFEUysyHbAgbaKyzaWy3N/oRnDCDIgZYkE4ue97YkB+GD4odb+KkZR
BZM+x9UgGo2GNYitMnyubmjJ9kPdii+7wlnT5T/aL3YHChgmS4c/CKbAv4lhAR5g
f6D29T3kUSjMLjtOkHjbe+/hcdLcZ+eslJK/1zhbQ6GqlKna44GDjuSMCTngd1Dh
iNXnXxRGTKeOo637Dwta+Zo2BodAMLcQAtnVQKbszDOHCPISdouZLg4BSnS4RpCa
fW4xiZ24WI9DGr/ifIRp15qnU7C68FccHQWy4c1Yex4f4fQNjpjnntOTywO9+jon
E2EZdqHmp0BXT4JbVUgTOkl4RMSJw/ASlEmu4zFt7qdTj07dzvTZ2+BvltkbDoJN
jYyAlRZt//UW8eStmHpcpHiI5nMP8eZuKPiQSvTraEbTvv7UkTqaNqjhXAValsbQ
LvTVHVW+ZU1a7B+YTNRVdIooaSfcEFu0gvHlN63H3+VDx7M9x54H6U6+rjV0Tycx
33IMxwBf8iMmFQ6tpHEN7ARIzzeTuEajSRaa6+4hydn3k3e2P0emvxNxjYmMxHo4
t1Q0d0/Ca8/T+cFp9A8ym15WVXCba8CCvtrbsNmDo58Ae+TmzHKbeOw4OtPiHkNi
Nk96kxt+2iO0KY6o7g1WCoIJs3W8dFfweZVgCG8ct27LuVAPl+ksQdeyzHYsQWq+
NhvvZ6JK8pkJL9U1Tik55u5rxMdV0WYYg1qy0dSMmS6BKaIPEsMpJQG3wborbBDI
VnrF5Au71THJ+7ufqkdXCd4EDLY+kisoeDv+0mpFC18bNREEdmHwYiM+RDUPl7rI
x0yFUQRQNDcQKc734uU9ZSjFYXj9frAVS6rVEjoO6F7pP6Jux2Tcr8G4mdA/36n0
uTH0pb0tDwiGi/xJazzevJRspHIeavsZDijePIiwaLkXgSqWhCfhGAmS1v6yxAhe
OKyDV02bZ4xQwT3QcN+2Lv5Q2uM5hT8lEgJfNIC52PZX+UOgufzo42TdBjNAAsbf
oeeQG8Qfw6Sk+oHML3Wnc8GIAhmxWNgVMOQBWJeyfJidQBlQGCKJo/0tG6ryIKbL
4UjkFwZLrXjZALlbK16kFgk9O50a1nkInAWlmSPG1K9eMs/zVPphxKapqY/7whO8
5jHiuBKYkQG4we6ao4XCJJH7fkWLD1S9iVs1U6x6OKddUHdvEqd5zEgYQAmlf41Z
D3zA5IMshLa6hkdaEQkJT0uw5qz2MCJ/CCMaqAxngzNL/xw3783lqcX4LaMMLfOu
Lw8lSkj2BQESSsSrTM2lPFjgY0zqd5SDLQTpByo99XvLEPgrIETbrx+pdR9ITEjH
u9pFEqdF+Al/9WB3r2sqvYuIK98eGG8q5CzOeUGanW/LU0bIoipUFwleKo9iDwki
3aPOxVzSN2WIGAPRDBtg5bWpMuucAACCflMorO0VPL6ct15Uye889qnN7TaAgKZr
2Wz5R2s89v11CsMe6BeliEypz7kVyas5ABdRNzRB9fi5AAd8fwd6OgTgdUvbbWkM
HZ86Z4LLsJGIidwUb8EXn039tT6R67m3/TjkUQ+44bfWtWDOdTcgnAek4HOL1f6f
hdcF45iRiNGHNfaAtUzeczP9sZz6KNmcgMOkExagcz2eSZhDEqdKkZ/3OfTzuEaj
IVONUANZvQA2YP8QAl5JNSL8q/QVWwLeKw/cmP9dmTnR7gobVtrKoNUmaVbXviYu
IKqAWMer8vgi8mcCrd8sODaPDwWLMJPp4MYeHXfbr+0h0qx7nZ0OPW7uwbdwsujh
SUUKmZ6Bc6JRaGeCyDY4HsiVRbqMmpz3rqTJZ9d82Qlt9HgcQHXH2z30KLuKOYrw
PeKkcIZggtlIsrgkU61cC0OKB/VDOeJkwsBYHC01xPOtcpVz5Q2unX0vOJjDYaGW
oEPbYCyvxbEwcen+dyt/fg9T440WZXaSHYFfy8hXN+pYlKdEClSVuSIl6AtDPdtj
pNXtFrXlHAoW5KYb+7lIFY1o3NirsXu5tpKW2YTIUbeLECFuiecaqmSShlLAfXJp
0RmD1XN0NgyYi499B0+CBosOL+eNCPrW0c2+YQaszUcCDrbmucNCHCc+h4a6rRnm
P4rPKG/uGbMW5iaCP9TtbE5gu88//Aoki1g73fNLlRtdHpPKoma0kiDgBqgjfEgv
aJgEKao08BiL7heL2kPEHvykzJiaj+Fc+W9lG6k8RoE6bhUE5lFvt4TwzM+p9m3d
FPqJhC7xb94TfOSELJp0bxEWfQeWHnHlIBIiAhNtdJ34ab7QaMqlygpRVILIwKdj
koZSlWJC4HnpbIqGNxmzpcUIZ4W8+Q+wb494P38OtT0yceWe5UEYcZZ4yH0Z9gP9
BE4THgOnAe5/Zr1mMvzH2JJyq793JcbHQVZmZM3Bx5WjPvZ+NX5b1WPn2XWPveSZ
wee6ImApWIEnr2ZQQvmE+q0o3jpma18HmkkQABO+I5AdxpyDbTup/LE8kbtjMqUT
lWGcIykxeuZoMWpNAqiyHSg4QDx2pwzc6n4RA2nKhLu4vqkXGPAVztGfVInQD5AB
/ojQ/NXrUpe37Ahpj9rMzQhc6yyBbalfb6/nGC4ZO549qoN/rgZT591MmxlVeNm6
wVBHSK+BMT94rNOmO7YJ7rTkyCu4ZmyHVYjgKRPqE3oRwKWbbu4nPBWeYrDOnxQV
i3O9lC9lWUGbe+SOs/EbkxVr+vAlr2dRf9m2BVIHqK26wde8FrsbL3m2nYFnXeaz
4c26aH57s5pMXMf7y9jvzWTe98bQuHV7uG0kWsri6CI0hAkN9dtPCpgmQGEDHVeW
AQWyT3FX2TRqa2oDg3Cjp0gCkC+23p9wQx+azb6lAvk/XfLphvWYyvScz+0LUoIl
8emO+ZX9ociiDJ45ZZu0saLVcLJDUY4eEazMauvNnVYyhK3LsOyOBdHWIwkJ/0HW
lLHVU5BPMbakZu4WEB/B30oxw4CwfVH4Vdc+zu1ZC6eoF7KIGi9HUWvi2o7ZsKX/
SAHJph9MIPtLoHchWQY5meT9JmAgM1De2ExgT48Kt75MaCegIjGcR2RA0ydEZ1fl
DKk6f80VYSSsdVNfXPMJ8A87Zg2W9sCSr9XS8kweMqWVt3G9i9T3e/K17R3jDQvF
LHFkkQcDximn3bZgiwHy3x6HuwdxoQr2M2Kmd4SiSSw3o5c1DCiDJCSMEoZe6Ua9
0Iar2/8cGnWmVLtxWl+IKHAv54Deub2c4IYxUe7ejN752CNAWhrM7f+bwAJict87
mlMQM8khCh20YPFEvFJFlxYYHrLz3Aa7um6KdMbtyXmyzaglFGGZx0k06WGHjgqh
QESN9G35/asOIgxj2AXA3FsxSKJRC95MPN3r6104sajV6+J1UYXtRK7TWsjGiQD0
JPhuSXu3uOJOjt7CHJX16kndkI+2WIROzpl8pPEEPI6n7o/tQEWGtovU77fpu5Hc
4Tl9SmjYVUv22Gj6dg+gKrxt1uu1Vb9mbe2b4wFUMdH/Suj952IKY7aHsYrB8+z3
rZ0D0osoe2fKydXpqWBy/lzqqVxK03KvKUvUaPFO9yoVlZOmi8Mh/m7I4GTh9KVz
ZCkp9v4PmNqrfx84m81ERSCqg6prcOUOm3hhS7+Oc/+HOAYemEIE41H4KIoK4Cgv
mbjY/KmzG+pRh/k8NSc6hUiTkx1Ft/e4n6dwDJtbvxEKl0mxp3vDR7/yHZRlGywk
jSX1dVSnlQNTuXvKlKtUiplLMZp+GPmDJIscsy2+FGs5+52Yd1t/aohCtPj2Qd8/
tZTTFlRQ5AUZBhT5XDEh//At0pfmtW60M0ZvG0HpivLXkxZFTLRT9EtXdOgeplKW
j2Q36LRvNSEO67Dmqd+HDokR7iBXHh/+X3m1HS3KNaUvkjkVxKRJfi6qCxSO6XAd
8H1xyd4SdXhH2IaTFMOwc1l+hlEcMM423CuyJGWa3KRef7VsBOJ5wvTAi05vQLwB
wJjpNSyssEjD8Nq76BIryz30aJSCJraGngKIQ5Pz5WLXHq/O3PNys7Zpi2Z63BaK
1op2rCsUu3bgapM7BNCzlk9XFAAe2yznpcBYGtU9401i2wNOVvW8+CJjwaBu66Ld
BH5VLpr26Ojy8ZIJh/i+5p4QJEREJ3k6xj1j1sZR7x73YCCQmUSQ/eX3J8nwt2xA
Tef/7TmC9ykfjm+E0A5FSLFU/2oQpfpvFv1O7sntWGYiUZADMRL7OakY67jW8DjW
Jzofs2zUB7lG4eHol7TaMl5N3uPNH64vsdwoskCYCbmK057HUFciSrjovnvekDNr
WXirGuCAa5V7MOui3TBoo9Hr/pClJM7j9Kda4DaJbfJbX21rRXxPPjLD04flHRIj
Hz3QHuc0TbiqTjdbzswtUq9+Xss0sajcg46Vk5XA0GRSrLJTxs5uStRGzKRqIZ8t
14Rm+kqFcX79iWd9fOSr8hrIa7caiWK/9dZLma8XrAmn3pBwdMraDyGJ9qY+XsXU
/MpBf5E2yPpDBV3FUbYXmh86TeysgeuEesVx/7ompiN+jdCcTEFkMxo6gvgPnV+J
ZtYDkyHwa+kl/FD6jzpZLJhRbl+wk+MA8ZuCgx1V0y4fAObeeYhjuN2FOKPOf9M8
Cg7Ms6mDlwxDuQMQLYCcbNTRt5IIvT0g35Mv270re72+R81T+wQv5fvxNsFjGOBL
BWdfQ0TwzPp78hCf0lv1xs+5XwzHgLmL15tJ39HDYBKX4EkSsbbCH3zzsGCaw1QN
FU4Sq4+03cj5/Dhmul7IS2TNyEINHisjdK6pbBneLOoj9qjz4GIEyv40N8HQgqnp
oCkxRN/6DA/Ml8y/p6exRsujO4BoqrbFXrd28Bk3Zn4yVSaoEIHqfHPhLRvW2n1X
qXAMkNAyb+pu1RZBP+FYi73v+MWJOIu21R5B7r3ujQ2bp5Wq3mPHrdzrJ5qP9oaL
uyEL/RiEaU/YE4QAhGayzWUDecE5IftD2lFbGhL6LgVSi8sMLORSaga7Ih8e8In8
l4/ru/oatYE9I1nmXqGI9F9YOQw3wncAXyQcX9HzRsJd4rFxLl4xFDNxjE+JKdlp
S2X46FISZnXyN8lYqwzudy4ZdV8bWnIsMklQJe1YZP2jidFfPqIUSmipipxcfphD
Fa3vb3NE4zPdtK6riLgXdwBG3ipQbQGb/HEZdxb4HC69l2A2ScvN+hiqnXX7lm+y
IxW1XyW4f7bhFtPFbNBQrKpg0NJ7Zmlj5JP2v6eadOLmI2GV9pTZK3zSSNFRHqLR
euQev3MzSTktvOpWgaXSdvIh+TpI/xeCkrHRRzUFJgxaR8L3EIHiNJouV8WLxYEN
+vK634NEx9/GYeur2DKGgyOyVkPN92JLknp1+0QDfwaQrDTsCu9MwUMgW5NJjteB
4G/8XaQispF8WP5Tb1SdwYJ7OslDg1ZzIt+sBrfrfBy1SvoE+Mzx86c21VLkm2eC
vQ1MDvZ373Sw219NiC59X5pVVtKVVzPkLi+89UvK8EUzx8BCuRO/T1ybK3YcMjYj
v5O1qHAtrZ348j6krY0D7tAQ/5QQYWksCxAXnU5pBpy9w33wj0NYGeX97yWNGUdJ
mfq8BYglyKfibz14oElL0amxBQngFX8FfgC1zANQ7gUmyUoG4ln73ErgQzCvdLxb
wdxdLsH65EAtDcUA66Fj2UZrt708NgaSic2pvi/SutmzDhghUleR436hhTfQsAAU
H8EWjolLt9pG789gTsQ8d5bfmONUub5+zrfpYr5t1eZyK7aKXIGrFtG+CfMEmcCs
pNuIeP4fcKoyAZiKNCgu5NFYpGYf5Rvi1jbODNHxQldA/lmJu1qFyCFcpCTj0bt0
IfiSVHUoSy2AusUABv2DFKzeoArVgVvq8FXffLc9td7akFOcotwn8zF+q1/mJz6q
c6cV8qiClWS7lBtfT/Z7tm8GYW59Z0Gz6LeJIpCs4Fn6Wywgyxixw0P8ZHKRIw3y
a+hFATumunCVu8AdRvWS4Gezv6hChle2PT5jgrD622gplv5ue1uLNaxTH8t7gNzF
VFFy8mlVw0m7+Ux2rvdnCIWPc0eqNLUbgBwLqyYgWNgTYpS9kp1sesAkAAUxtDEt
6x7zLVUxusDZ/ZBPrekT4fImjYjPX87HHkaNCNR85/TYujWXaSKL02kEnfji7WYS
cdyQYknovSWnkfchfNFxYsJaH3xNguOWNN2Lzr4YzTFx2x/cae010x4Ed5Gv2Kvw
Vbqe8qEoFx2OUemBXjnqH0KjKBZbuqxgix06FE2N74i3n4PPuBGB72wanpxKRdDS
RSuQxjsLam4pSuictKbHTi3vibdjlV/tTFblZCzBISQmmN8HB590YvKLKk5K7K/O
wNoeC/KGAYtgK14wojnzQfCqKTSwgqrwDj90krdTejHhB/bWoRb77KIKnvRkpNew
Z/xizdXAj01LrOjdlBc9rxTyqsy4/1aQpE7ldJdRq9c71AyVehebAmG8fmGRfuIZ
HzW7KqCQZ7YO2n7vS6/+EzCtJXXKJufnateTLGAcXJONewqYCtQgI8NFulIabuVN
PEnOkeaIQS/JcYSdx2pyou24gpTV/TeiYHdlkJeGjTpu1YVuaNIGteCARbrQ/kBx
e8ji4Ax7pusCCO4YrBfgwEjCbqQgjCSlZ2jyFkxNbojpP8kQIr8LBWVUdizbBel2
bmrw5idm6y7VXO8hjv+6x8ySIn/YTycl3Qe7PfO8BoAtptwzyqHkKw6d6h7cvFRN
M5kEWFqowfFzIdt5J9ZS7fgQi1MVC1N/9q7XfdqeOHdEZGcD9slIXDzoI0tb+700
catmZchLM65CH0vQkTY8lidCXW/SSqz/gtLrf9cD2sUKEbD0XcFspecQXF0l7cNU
ntFek1+Voup9vZOuFTi8SzvOXmtxgdmXG+bwLYiLbjeoBV9W2bNzRVWWuP1iBPxh
TA8lCX7hwPnVOJyJltFMeyV7lQZevRLkEi3PwvE+iVB6gmbZJ1UWp3/xiD6cMHEa
DSWrYGlrWvZMk4erKogYEbwNI/iuALgi8ONbmaKIZDD7uHTDTadU0vEHyrRchWZd
x+SkhplYPbARz2+MQLNZWBd2RTA2U7cFFHjScEBNMFuGBQNioK7Oo1C7yGE6pHcX
HXZpx0UucMwdrqp77vCbaeIh61EZVD3sndSDeSQuEMHDECl14XWQ1B8DS3IXKcPk
RLOl/xFz1DmPDidByTr4TEXAwLxeXP8Io+9spxogmrhGJjnX+r90iXJF11BTSuja
uIvkv3X0rXSsXH9JW+16s8aaosfIuK3XwxOtcqzqLJEUZSdLu9WnSWSI22jGrWuP
zuuI+FL15Vw49iVjXbf3S4j7R0b94DZivQBrdzQohiaeTYByQbbxb82IGxM1DSx9
ll2n44CXYpmVapomDHjINcQDGwO93vNy2wVXtF5wFnHIXoWEEqeoEBQCN5CP4Fz0
MbuFqpIa4E7KyClXIS8aWbqZftqQZIVs9umyi+G6K+OvLoKndBDlYRXTGEfbrFR3
ubK3U2tFTrHZF3F4YWel3nJ6LK3Z2R5gSDBLq2EtULdIRSx/iGOOh4beQcHywY2O
QkmYASDeNVDpMLMt6dVrYH5B+SgUuheY8IuMvX4wlGKEU7KtsuZoPFKpx3YmYNpu
N4DZtwGZ0owGIln4XgRU0bdCMOrandWFGZUobrM/1GB+D7eVvQXPdSzkKnFZX+Ot
d2zNr2P/8ZDZMOXJQlvg7ruZ+ae6FNeUHXQrhdxhGzvmo5ooDVlUw8LcaOa+N1IN
1IDXmvLPnEhhq18oevDBNlC38ym1R+zKVFcQnFKm0swsQBfhXhiGuPZ+qXJXYZm+
7nW52nQeY2RUakr1Hn50DKJtCZ1CvJGxVndQHFfkOsDEB+KzwEjpOmkI+PlTTNw4
7xv278Jy0pftM1NmQnbkF+M5zQ+MKQF94s31VCuhwF5STf2fUvb0baMzQLskj5ll
nbl2jyJqTm/Z22NRFTIkKd99UqkfTGZp7TwpxN+ZcjzERe9q8URX/IA/oYEOe9Xz
HWzCOAkM3NKLfAun+QzzRVG2PP+1g1gv/KbKjcyoP7oJE7GPxK6v+OnWz+U8+sAP
5i8+JRjItqXshb4oAbUE1We7k9WRbkV9cpF7aVPODd88qlT6b/jwofuYIng345wX
LpCxaAgvXtoNQwAVQNdZZzdWWsT7FPWKWA7mXUHW2FykYFECximjTKV6TyyQ2MR8
XS2HchW4xGnMQeM9BqNaM5pLFOMlxIBAciWh/9LTJLIu2PFXy+yLJMAFOd2QeWpo
xCMtHZ2ehKmbF0H8F9avTRCtDEMkg26I6tnSVRuFnrIw7ja9/ha/amMbojWMiqeF
W+EnL92yqONG/tmRaRk64g1gHN4K2cd7OeImPO1UFExF6r+ZfduUb04PdfBNya5o
hN3TjdZQOta36PgA8AcyxRIOf3zocCZWISVeTds9NH8dcc9vdm52fldxClcdcgpc
tq3Vge8o+U2/7RUh9g2cjjC8HEQBlEMwjMzLCVFdlCIROetW1FBm/Hekl4tFLyoY
hZCPvr0sD57ocaPV8cYQ5AImNzxDB7VPJeqBUliVl7n68NCZ+yasE20X91jij7Mk
irwaHrODKjj8zrMTW/dk0gT7s9n32Zc0OaaJqppgmL3AfsiT/2XZnBk6SSjqO40J
G5N1E/mFXSr83YNh9rdkuWSMfGthQvVQvNh/tZrH3PTIYhbvEby5tKMQs5LiYtl0
vtnzRCmiaWLhPtBKIsuo6cxKnpkExm0Xf+SYObbVf0w+YwpghoBBXiGY/9j4DYbh
19hMDNcafkfprj+cBqRgPvyNE+yn9l4lzGQ9SDtKRANX35twv70vCkbRYvIHG0KZ
1EM7r6e7TC+iZrjPamYk+d9b41oN1JCDVnKuW08YFLModhf1qbibEi9QTNfAAKT2
/CEZCRkT0YCE8U0Iw6d35Rzy90tdNs2HYT+vZYko/Dd+UusizsGKuiVtWQo/6cWj
mxLBOXDbSzjptqcmxi3A2uDAZYAxGzoOY4tfs0nsq+ihM3teovzlvBqxdbYzcxmZ
4eTxn1D9859+doCdlJYANgPX+k0Qclke9zIhYmAseuOUu78i2Z8wXYzWgN1jih0n
s/3F29o0ReKsQdT8tPVSyAYBs8PKTELjEq7A1fOdCxhgEBu3u72Gjd0ojafe/qPg
IvrnG8AW8CplfokPehRgxC+H+gNTbQ7IAizVrpgnVGxpfui1CMuiokcC1IC+eKly
cx0I6UFQfgkAJMoIInqumjLzJWLMZlwF4PTO9Fzuadk2uEZcsS+qUGIeUdk/22wd
bRIh8XSCz86UadojLKwAUpPTEdsZIumX28yXyVAGBbo0Llk8Lt+j1Ho3uv27pVWj
yRuTrPO6mBQ1QELWdOAU7mv29HrkTa0f0Ch6f7b1sgbQChBxidXudOn9NMWT+Ln8
GCxkQ0aFG30dhL8hNCCqqHSCOO00E8Fk3H1pjyfeKyKAMt+90B+nJPDiiBMMUeUQ
GNOsejXOVR+pMJri2KqPb/jbB39Nt/lgA7tbSoETo7BdsnSp8+Bqy5Sr+Tmg4Zph
CabiHURF0FrM1yRa0fbdYl3OjwoEr8VkmsZNIIodb4n828dXwMeCjPQNg8kQbzCo
WPqIwuwvpJFJweH+L7e83z6LFVfl0kHaBv25lDCllTWTHAsyFcm+t0AooCy7rEQz
eACRwKIy/85rdHiljPy+oyYPLiI2GaMSvFzTOO8imAJQSSAgMGDHpnviYibmEz/e
SV0YDeeNAYsDxwdBnU+QZrXkHj9cFJT4ToMDPNcQBZ8cmq0qgBccnPSJ7s6QCUsZ
thyFugvwdn1ScJXCJC8qRg7J4Z6sc7nmnCT6mslwMz+HW0rDGBc5ke7vbbyssFXd
NYklcy15PiQZi0OmAKTwt3C8hrnu+X04JhYz9MkFO3ZSuZypH/obX3fNXJuQp4hZ
srkRgEmcC6tCfWzflMLdrhysxobPFi4gxTQN2+1qvGJa7lT7Wzjfo4MWYdJ/GcuI
8w5ih7xqZ4sOM3VJSPErdn7UmkR/Tvc5prAELFmAoU+D+QZ4ZRGxWyfnXkxocxPp
twkAVHkLrvuO4A+QXqdXTXAmJYlYjl5L/WbUMRxvj3ipxff2qylZ4a11TYkAuliS
137BrtMo0qEiL7XZIYuyo+ONE7cJCD6u42irppTjT8VhBCDVeoyo1g7nP16Swe9B
F+hP41OeapoqAYWrADwlTLMWf3q7p6eEgEs5394GhvJD8s7ff3NeaTi0zJhz52vA
nQsPlETCfGZkamjGduy45pkTHzUCtsv5VdBtYmKz7uptNcCzqGyEBMW0727fBx6b
GYVha4FXaCloOweecaDI05oDV1esD/Co0E8qKphMxbPc5kwEEcTLlK9Yb9eH2ZsM
uNSSrQMM/W5hpVQDtqb/fy+2iciRyOHqWNsWy3bJeHIk5zUiyqTN6QuYS1E7jrRk
v1l2Qf29sjuqYn+hPZlN51o6o/HaNsP7ND/ZO5d8tLP2c1KSahF7pLHcCOOU2QhY
xRrvdpIyNZiG9/1BoUtcFJSBRE+Ai7eO8ESiq0E7+wbp9cWpHjct93+m1NNluXWx
BaFF9EWkOFdIVyEWiHe9vzOTXLpKf98dGEhr3/whcrlnt3Zz9ONkcmHnzcek2Dul
cBDLU2FHWaz4wCVXpx3OL9jy1oNCaCEHtFcG09Qt1BP3Oia4TA6kidyw2zLPBdXm
l94ubR4mfdjuE9rqkGOQVlOMgbr81CCyH8ySIupj3vwxPBstENcCGVjaN3DRlDug
pDVmtX0le2dGFfcvNKyd/J9D/D82BfYWg1ViTCijpb2//4+gQoXzoWN0NqAlzHkS
KEXRNLfU8M2jcMpQfJTuZy1ZLlInDY3rANivsBWf/llxGPetpNSX88a8F+SkVc4u
DfXYthugaBtVllVgOYUhhkJ+IuXJyRAZYEB2kRfqz5cd0yMp3yldLxw+E4+4M20d
CvELLxNP6lWrkpG/4HYD/+zBks6R/H7CMbET7dxiufFMkAYIEJnqDm0xZueI0ji2
13Ptw+IZoh6kyenVGdbaualUJ+JjodovIuOcsTLMCl6C/WTGPfIQ2A8hwqyvJmbR
QbjJdAVd7Ap4tjN67cAWqRkTLl0tbZ3azI6A0HZW/Zgsil5oBqk2H1dOqsD+3rLi
mrlWVbuQFfgNb8NtyXqkDJZ5B6dF8nULr/YhDLRnVZWNom9FlfkO+bwL/6AjT+4q
MvpU6JMl3m5dobAJ+GmdoXmO+cFli4B67PqLSWfCTgdfoMZla70o8wVK3EU1rjLM
w0VhCk0PiD6Z6Z+7rWpGW/hagBbxhjWGhEkq2gu7y3YGGDflA8BpDHtciXnb1fzA
T/fsARR77SLzLzilZvEJ8jf4wpchdRTJy01EA9qq5byJfr7AhXGWBTfl5rszKsuS
jOdarlUpTWeeZGtdozVRndrCxpyksl0ofg9xpzLwNZHOo9ZidZPzdcuz8eQ0GDOv
A91nYi8PvhjtchG1QEg4eEFXgnrBYQCEEccg3yQQnfeGRvR5a6QhzIfR1zwMoijm
6aCRpqTY+d/nbgpzFsM1L60iXm3lGb+Pw9uDz2qvqXsaplUbAWSyfMb1dmUyTh76
r2QLIek6MC0jJv6WDP4i8G1lJkTMzi9anyyRYiFovghALl9ay0h2O+ma/Rt+0c3d
P2v3HGMKyLGZRTjXH3gpUl7Es7e+oMg7qqo+MwuziwPdG4SLywNdBQpL/M9hQZsr
ZfIr2n0eEqSU/WShnSOHthcO3oh5A0SpiwZ2R+iIvLD7b6UeSVDe9kfYnDOfu9QA
y06G6Xdc8Q2HiBGRyN65+6Q8aDQ5QuJMlAkQoFO20SWm/aLj/hZKfB+Qrh0ImkHa
FtSHyZBsDGDFMzQVJXVlNMXMABTRLa+bC1oFXFrljV9LE1DWkle7BuxiYphpMOOo
DiTlbgVbiUV5+lRW039GwDUxM2rcbIw1eAg8Z67NDMfLWvHasXIhRoiIjnqtqVua
A1B9mwBdy6+bamVQZOEz9pWubcfUe+1Aor7dMnVLig+7Hb0g17YEXtHa4Oiv5Pkb
o8R8AsFO9yn5/Ojlm2Xl3OlFxM31sf7DTiSJFDsKhu8gXZJkRZ3d2ktNjmjrs9pn
1ijCNema7WEcY9OFQuZo36kCN+62z5D+TCsp4jLJasWWlFDHxmlzszLddOp43RLw
L2K54boLSHUXe93gQLhTMKympNbg0zme1VCHyJ7UfxQymmVPkok4R4LMR8+KlTTh
FbGg07rscM9iwJsaqErBHVrsHRI7xbW3DB/jThS6nvvx5xcskq4vKhOjHjiPFO/R
95MWQxey62rksU9Bi9DkqomtQ3Umb4DJiTdmrw+q4hK3YoZc+Kpzb2fXmSOQQWwc
GiMkww51eoUcNXNcwGyfuU0BiYCpDi7VxfYHsCDi/B66yMQYvj0zKD9xP9cSc42d
MVVFc9zV5tl5PaSPEjf9ZKQpZNg9yBi0ZcCZCPrZ9BOU3UiQo1/Hhzfj+Ca8t6eq
JRoXN1segRvC/GEeheff4jXhUWH4DlN/pboqkK/gSxxzFxcrNnLOT3ichcnECM9M
mSMQy6dDC1DRn9agiEOvpqiW5/BD6jWaX+ubDCDev3hVE3wiuyYnMSMI87JSmBD5
yuvtldc0s4xibcNyW+Z5QiTjyaPXj951b1CLTznvUloLv7uQ144i+q47d4Mla2o/
1/IGWTP8lIfrVebAYolv09uGZ2LPuzyHBxBegxcuww8lL5O8y32AgeqSEeg5UCG5
Il004/3PMRzxY78SsWjwSGWmOCL9sgyCC9LAIdPtHvoAXkdkb9q2hk/vMv6G355s
q9izE8oGxi6gbxPR/rjM7UYGLRCoZRsCdpqUU8W/vcWXWXv+7xzF7MplYowNf9wf
N/0IWX1Ub9AyZWqeLbeBM3e9Ccb85Qy7a1zyNhhAlomeLHBmUVNuACZwwsEzHEbo
h1ZtGX6GhpYkDovUMQPjB64dEMn8csR7lKhv8kDL/UqZL3PhO4g2eXqo3BsTQxeY
N6jokXY2tDKxAfvKr9445mTG01w9IxiKOnOzxTt0GfkgFPOGWqg+SR+xute5Avt/
9d6mVKS1Yje21MX39Qg+KvXLYTtCvlBBH1MNIvJ/pDqBfotaDLPsyy+mCaUyDnGa
2Na+wGpW4BatAShbhv3YwARRYtN8rtq9wpK9Qk11bq5ia3HcD9KE3iEQLcVtca3G
py6e0ugnShP4PzUAGMScXSEf4HJQkiemd1r/UejaXkQn8IixC0rpt7TU5PkNKLIs
k0D3eqVonGr3YmRPw/OcnRd13p02bWBdrC6/2ZfbK4XqlFbEYobsmuYCiKW36lJm
iGDE4yOOl41X1rcEtWIm83Tfnd2TZ/strgs9pTso7hrP87oL9Peh/pzN3T18FDNj
2MameGylCbKiLJbcAhyTThGJlpRlJS2avkMG9A17auTRSjuq+PmRW0ZlfwEA7kOG
FfqALCcZSEwZBlVMIpR9jzlVcjuohMoMIF9Y1sEl76imFVFD2lttWqLi+8l8Fo/+
5EeX/wLtR5YyIw4wzwj5TlRKifc+SU2/dJLvq8HOa5Zn62OgOohDjCmBpIusqfog
JJo08ZheVP86SYm39rgqm+qNdcIXTNfxB6uh3hrsYlrZm01IKIpRhSNZtYSwJqL/
s4hf+InmGw2r8pChTSzNBUfhCLgcUVqe4hBIfjBY7/N8+tXoC4P1Vm6amonGRHbS
uluk93XNNE16DL72TVf9ObTZh8dCpJwwhNhV9uiIcYQjEyC8iMx1zdXls2Uvh28n
+KPvd9uAmOpESr3cdyYSvvI8WghMrXmNI0MULJdDHIh9+ZFM4nz8kj2SIbQkUHB+
nqAooWrxo0KX9y0GiDiTXEK3B8UXXcCbs78nCeT77i4hVsY1hfxCvbErGChUk8cu
4cG2tCwIGYPzA2LFLZZrCLhHoZuIBRFWW/KQ8wOBoP5/eHytpnJ8cRFSJrkHlHbJ
rDnZAH7k1o0tqM+pzFaVVBLa+kX2IJT+TthlDMHw+F0+EgbbroSlwA4v7pGFnB0Z
8JhQhbAVRzWpjR+cS5+aTMMiFnGb+hey2zIEP5+DoT6F0fjc2qQR2QdKdD57GOPI
fKjOTqhuC61Fd58uTEZc1Zwr0snmAiJjeXrkk7qyekcKYyLHPDVmibUn9bMHSEUR
FUsasbosAP9QTrFA27l7zhOcqEY99cx15QruYe7XPAD6rusoRHbMIdSgAGbXmuee
sxmqlTg/bcqpIdApcEur4fSVXi3Hy2tlY+UfgiKbZbM/LJReg/S1hvmNlkmf+5bK
7QqD+2ra3mILbzdnRMLE19SUlEiqwf9iWAoUnzwfG0P5GSByFsVB8OYX9ze0/Cq3
c26jvY+3n6GuhoA+g8Cvg5Xt6aweuLbAEFJUn/jF2u7ZQm4QAbBvGOBmTwLSGG+s
wAgGfG0W+/ZS9Z0h0xYmPdFju/FCLct0is8NziaLQGd2cMLF3/VLrJn3IyKk37xu
6xmYzCfqZnxc4HmJAqISqecs87dkTSZoh8AKGPOnVhE4d0djuyOxOSjeKKjtdZFI
XytR+dlDknMr/WKrRoeW71VYLGuTYprpY1oWS9mnpxdJf65bsm6MRO1Um+zqAsXv
eQW5P2EKmvbJcyk1fImQ58F+FAK0VQdqwgeGEkqlb1fh6aFPpjAHrFfsiw76Rc1q
mm04cafKQDi7Slvc6mZ1ZLgShVU4wNN/Ltum8R7oZssUv9uxl4ktclFrt6OFNsJX
K5N6fAygb+ekLJhU0Y8fG05ht5Q4Co6brNV44CdxSLiGrNRyQbxrCbHVnq9cBoaZ
+mCjmGMYOVprMJvMuTBJfo1p5AsfGZGHn3gf+xaH8v1XD3odx4XXQxB4bFuykdXZ
rcGLqNue3h0gc6ttAkq3wTE/3YfPpaGZ4rP4uh8hxWMlBhUE4NiUofwRwfzCYq8A
sD/7FpuhYXZNbAT1zIKdlq3yYJ+XH8keaKzXiwsW47/Rpic1qb1UHOSaklLFijfs
7VKC3CIlJ1uWYi+AvwKDXP9S6xLyjhiIrJNF7K7YgBWLKOBd+R+2mSevdNifJ36M
lOgqyzM6Cx24zUx7ZQlerk/rL/lcHEr//H7xZ7Z1cfPrH+hcReUlVngtFEoofFli
rxolaiqMheNiR+qOammbgoXqwpmqqm62rZBhFJs6CEqIkAJTcZm3noQxgSXskWo5
WOOdZwG4t0UKigruVUC3LKvOWxH2Bet4YnWJdMeA0Tv+kXDlrPG8CsKJ6JwtbIcI
TpdQGQ8KGJWWVqD/C7VpA1jjDtpYOcarUMKgR1TGijkr2NJQEZDZPxqQ3+OEAZsq
wOF/aSWQ1U+NjgFJIwCb0fZGhan1gWc19RvASBuJFnc7CK6KM5ZDqQB37Hytkblx
TbrYqCLZffW1YWRcCeCk6aYCie00pCTHp6d3khubAzwJjnRm85Gd2BHUJ1Xco6P0
ZM1v6TWHCgVJ8v/cWjcafaVlG3NZNS/oP8B7S+z6Fmrvo+EJthHFP+tcrImzV71D
171Nx+KAKu9AEutu/axUV1+n3Mxr7bd51tQnPnvesxdn6p8VjOVCkY2Hyj8tnUo3
9fJhktVYp3R8SX22Z/Je62oo2c9bfd7fGJzZH3WQoSDnlGMDRgQ9i78b5bP/fVgK
8gNg3OI1AXNyDLu+u6YBhc9XNTN0aP91JeREE4qedLukrpdR/CwCWMeHWWhp3AMS
fcZwb5zJxOPzDcpTQRzX6m6TzusX0MDraX1pAUIFGnP1H3taCR9wA8WKgr2z5Mht
J5s7MWIYzkERJXpoyKsUcJQzVepVTBYmJ1U8c5D0quiE+4ENH0E5yZdbFVVyVRtq
wLVf6KBMAgpIc1TfwrZWCkKeCAS/U2U/JCsyc33GEB6ZsA/gyiUZdhSzMJ3LSHBZ
VwQSwxH2Jviy8jG329KncWu+/yDSlqRoZNDcRmQHavDILipGv09ssO/oj5wHxsAM
4epMZT2KL0mnYlnI1MLWwvSmpoDz4KWVC7dS5+sgRolD4qFvMJkVwIWKUp76NsSm
5rU3BV4bYvDcDdPuCOgQOsZiLA4BFEVX/Qu4MgBFqELfod+hKp4YP92m9fwnM3HY
QJMih379F3/0EyP9h4PP1zQdOAADtAbFmVzOWlh1gYrWBNvMMhdwhjNOfsD6i8tI
yXAjTzCfpMLseA6G6hJn+kZR0jCmP87FpEH98ihzNlFLV6MN2eV7vKHZCw60F9Yn
zWrTZiAN48rIBKneRNMHRkiHy5xXkWnZnXmVnZtSBtrl2AAuuTKUIvNxi3cz1rJL
ieztrzDF6WkZYtofd8j6ge/Xz/RI+erItYX+UiVSFJlMEy9gc/emukFhZoXBS+X8
zl3abvt7K9UhIDqJ10BZdvv4sox/V+mSr0XPbwJB5iD8aDLXMrc7nkK0GajuTfQY
iT4mm+qEIjBDH8JFPuL/+XTWbNe9ABvF9b6nXl+nnS3vMXUsvD42TZfwKhlxRebJ
N1Vu6+koyIHXYWVsDQ7yAmOEbriiABUIgFFGJOu3gCmlacvTL6LWvekt1eumxE/B
lM7y5w4TEHQl2tF8B+evNLoume4AJF+bw6nvu3czCg6fZpmBddd+5RQ7QL19vUX+
lPYt1iaiaU6VbNTDC9eGsPC0EOfKJnzjvoAAmqf6l4j0fiSdC6tXJtqSau6mAsZW
8yFCuy5YqWh+w02v+94t8LxL3ByrXdyRQX7/OWOje+qt2tLcLYilDvP+FIWnTGMl
EJyWsEs/wgngaCwp4IqAyeu7xoucKfq2RLY78wHg1pzyhx7QsktLwvKwobG2pFEB
PHrfZqR1Kfb9lqvhwxQbauQIMIl8sFwd5AGAz3MQ33FyUa1IVtJuQRor/cWX27HN
LYtMSZhzCUDgAoBNvyegXqZOXoUsgcCKz/BGRZcLw6+NA8++rcnsSlQDVaY38mLp
cG3xEKT/xOlp47a+aRRzr+PuNnXPb6cgXHqyJbFaXq/uUp99gh2Ci5QpoP+43w1X
rVGsu9UgmshlkpRpZhQjiRe8hB3tpqEpIYzgrPL4bnhEbOcuazsdY0ZxdthpL6ZP
o/b907fPIgcDnrOrxoXUxesYK+y3BYH4Ru1k9qpsNmATzQtzZYz/hTBkz9cbiH4I
p6fmU6RNjS30wwIRVplAdx8q79fAwOKWpmoJ2HJ0WWgcHYo5iANXFqUvRfO/Whd/
pPbVum74CuKCcFm5hJ1zI4PxX0E8Y5Rqv+EZ+lPgMncx9VaQCQVaexRuS7PXScRx
juj/+HivhGxT70khsGw7N/vfdyDgEbkrX7gM9d7zFZTdNCvL+JOR0IoZ6XN9ISwF
8SEWfSksfUgDhD6TG6sM+b/FaCQ2IP2WRtYeMT0bapM1NlD/011bFmQB6zouKo04
9wWgIFhSSdAgPFTxw6XNrqLMRfqJrhsagbVh+hCX1c4Sml+niE2LLlMGinIS5Mh4
7pKJ3Yt6abzF9PRoVrjxjYPcnIobEnNbsBmpBiUruXJzZx+lhwq+8pwE+5NmnkR8
vB7IClKGAcCutWUY+Ohebqh9E8MSKztse9vXp+pZIdzvgu9w0pU+tYuNvtzE60IC
3A6NNb+gG7jzhdT6ohvH5xdequ79J6ajke/8kvmL5Q/ZmMOxPzar4+6A0JpfZT7M
WxlB6IEzTLIcmY1Rq9fAq8uVQLTVdnFOCt3xsTxNLhZ7aG6mThMCNGk9JlXXJFaC
yev1X+erAayH0nHGFq+5t4sSQN9vMTbyzf9qnhazU7pTaOq8T9oz1sOpzx073Tjn
LqKvsRyVoTXzagn7ihHyjiEF8xZ1wqC96t4nK72Rr9Nw69HdZXjQGCOpdul1MtKE
uza+FhaPeOGkmdt+03dDXz/ySDG2/U/ag2B+RdpFHd7IA4bvjOBzRjxH/zy22qLN
2bRhlvdhKItbJrRFJoaL4vrSq5XGuKC6Z74XsjvXkp2ktDBMw1LmRK5+1bH446Qf
4hBwLwDfQkQBQ8x4DKwC1T5dcOjbk9oV/TfTcaZxWJrLPLo7SvdyqnwDz/lT7dQ2
se+bEmo5tco8+toiHj1uYMmXyIBttz/5GS9hkvoTUqbLuiIJWuhRCv/s35mCtr4N
VpmClWAmek/ErOx41Xh9PtRMpRJC43oiw0GE1m5IOoINZR8pJS04eWyif/3rUOr7
kkR1v4WEKUPKTcu4ZZYVdJIHm7ur9n27U4VYGVBkBB/kJXp3TTE8BN+dVqKICWnL
fHLaAWRLdriNU0MEVecFNvIowkYTCvU0UKwJciJaaEUR6VkDPckdzwj9SSbbu3Vu
HXLs1RFigl+V1zEhAGmYphcbph2e52vx1lPSUcbYTKou9BAIxbxD+MQ0mMdu1K2K
fY2gpboRkvBECvCBI4m+3eS8MFBxvQU/s4+MkjC8fMOCWCmWVK6qwdcf5b+C/yMb
aksh5El8ZSTmDL3okWiZ1K7lhDMFoJ7+0xnhYtRGHouhR3McvW5q4dSukq5Y1gKo
n5JbNjTQDFf1DuWuczjc/yeLuQsutrGOJsnwKBXMG/fZ7m2LyF5JUAludUQ0Qyfi
RXVDlMgPQ1fTXMtiqyHCu4eOJiV3k5gC8O3PiBu5Ke08grFKqX5FgSWXdpNg6j1j
40kKdPfbfCr6qd2Z4B2LWancmog8Thl255W0qMLMq9xPoyWMx7m/qtTqeW78xCJq
DCWUXe7HS+0HTqX+vwz2/1YMYXArTyRdZdRjk0AEdyRjKt6TTdeS0573ddajImqF
yfWMXXsquvqQEuZDndtAuzTS+BcEu0Wpafhzv498pCZ8npl7qTNS6XSiatcjhZdR
ln57ftTFuEJiOLWjjmlnl3rjXIJi+m/PSy91hdaNdfXeygotCZy/nQWk6lMh2VyJ
ernSmqzN6kXY7NVnaUBxZ98n4qcjMJSfFvKUHiu7Cze8JS+YdQIGQbNQh8pR+AlG
pzRlRK//evNicNgPE4pCIFb/55fB0rCG8l8S07dGJP0LjRX9fQeJxT6AWh8qOBwG
vgK5NLO7d78MHFNx09blxvH7xLbdqTIN/bVw/rfuX4MmXi3NJRZssdPoBdAo/Uow
ioHnftRjN36oSXv96zwliXEP+dfNLzUd49qP8XgLzKeyqQ665D0fijspcvsQsDf+
AKxILmhvZpUhH2v8jawTiuS/kkTT9IHeg8l/02bL8742ZfLY0682cqmaHmcyytzm
PoS9m2W8OCGLX3AZRGTG74x1bUH8/Ca4Jax88elqrCSlIGrR4XmaEPTUC6JyB8uW
lYPCCOkTOg27W9tAWx/bESVPgxN8eKQMcC8hH9/D3bJ5Lo5Dk6SJaq9aU5AHKtTD
Z+eFDWBBoGm4N6GedBk1nS3dG1zd1j2HXkQHn4V4hpJBBykRkZ1f+UQJhso/UnX1
GHkz3LvLkk89oz2M65cZmxD7L1hI/uHNOoOastNO/ZgLO5cOZ4wnmzhSaN3NvT7j
ucdJCx05Vpn4YAvz/9qYw23hjh13AmU507YPel0ACZ4C2MLyTcfE0osCX6zauDdh
vGEduR5RlsKxEV3MQXpo3I2j5B3XA9PiKhElNmsK84i/qZPZ5nSc3JB2esAmpADF
39PrprPpDVh5nmjynH5g70X7hkyDJMgSMmeJL/PSq/aZTryvPFh8a4s775fH+II4
XEbuJ9RDix8gGZSuPDcjDHL6k/YeOIuFM2rTtvMiFN/tnH+DBEf6FzoZFYBT9QhH
X069qS8Ldgkd7dWQJII1sNF/DTirKXs92o/qlICrL0MNZnu1WV8nkgQtTpV39Jaa
In65YowbXq6DLbRDXTopXzSQzmOHCbk+X1jU8jlAHrm2xwoyIBUvkxu1zbmSESwa
ZLqcC9cNtcXZ0/5utMUZqWB+MXLiZUy+139dSFp+CO8TVl1nCxsKcjhzVWKGKwxp
Qrb6IwJAVQYdI56d801wtDnk0+NQ2o5dnzd4Aufy0uUBJgjwaqsMsdf+mTH6bnS3
JRxuXvudeS2wqxyI+QOIXX/6U2pi6d4AVXOhWDOC64PdhkIeLXVCvKjlzP8lBi4F
aeEOK+gUMrzfkJy36m0eoRL6NNmGT6vgvp3koBH59JQFLDthG/BSBOUDNDPYVg1u
audg0/DVtywBS1FX3SSMM2U0FUu1uxyt6sa2CuE2rka7IjCBHcqPqqUL/UShXJ98
xwpXgIXOzcTSPzzcPrZuBTFIoJvdpiUC0MqbpP49V/qDnfh1B7sYfRiygTRQiiCj
12+JJ9/5eS/a9McbDBvBuEL3oQHQoVS4CYiHPNAcmLjPMhdV6o8VFah5AZi/3dDQ
9Ix4xzwtKYsPjXaNMW9+einvh0yzZoqzj60f/mRN1QsqTJKA9d6RJbqR9NSQUhAF
VctT49jkwyfx4eWuWqlOneizSSLei2pyr5yPaFsNeosOXhzSAZAAQQn5P5SHT6xX
4NPU+dc5nf/0TgOfVU9DpVWtF//HD1mAFVSl/Ypp0CR0SeQ66Tqab879OV/vgqL+
1FShJIem/VzQ/054bmnORR1lPS934A1tgeecDPfVZcBTsQGd6XGuH/XoXyCfCJ4x
JsGhMeJ6lsDtAeyBqZxz7FUd5LTfOZ6DoNvhPfPn6TeOOQZ3GDXmdx3ywWfYHBec
sq8spgtC4fh5rKCZZ+yhjrb0e+LJhSMvbuLi+VGAdjQbNi4MkPb8gwDjs6meNG8k
mT3Ys0rzgCMwQqGyA+8dKIUhof4QsxBdz8T4yVJfPFQUw7Y53u7laixV652cH6eX
B3z5H7OZ2aE5+2hOzcgQ79dVZrQDhnWNd4SCadNNsjJs3bL4D85sRP1k6gGsiOXp
iXv65H1Xdu1cZFOh1rL2bPgobj5Xh0PjrGM0g890E/xMJ7ekonF5LUPQmzi9ifMv
m3fUEtpIubsaQ5ViWrcJPV1e901ad5gLJvNt/LmU5IKCMZbl08N9TCp0snhZMlU3
eqTq0LEqd4mmlbzB2HC7PSqaPRnJatArrvDDfNoWGyydh3rylrGSMOEgnVplSrcB
zmIuhNQ0gWeCwuvunqiBTvPJCXFI33bSeLL3PgoXl8nHaw9NNQDYgaAukf1vUuQb
3aXH2qeZZe7rQcRQBx8EvOXcFxdwn6dWFskUq72rcYETIQ7IaFedfk/WT1YDpwzC
mpgNhFWb2W4DDwqdMLfXsytoqsqOZ3mMuo+YLGqdwcpx2qMFFszaYDtCikZh98D2
5ximG/rjMPUq/cZgyWgxDK2vzXQhzXvG123rJ6tyo8wxsIxx44FMHLOP+E5ig8Lh
ReKaUi99NE9TU1K2+3a39wZjDosQVBm1WVanG/320lgLT1Jmli4KdXZ0XkrpltcU
ALYsn3ryHKn5gPCdXwZne/lzfCdBfGmqml5TG5bFY1r96aCTrvJMb4pZYmqfmhKx
6s7pHpmUPDNiESDeIhLR9i4HPVjCsmV5uvFdYT/Iap3CAY0Z0O5PP8qNpBhFcT/c
c/ulxms9qU+XBCzFBBOeAJXe4Cb6jL1wAWXlmA7EHQHHCfQd04q0u/u8tJeSZ51r
UkPGUuEFlTwhtuHpCSX6+HdnQRTOB3QsB7V+DYBPYTZbf6hDxjpAIHoBDaL2W7PC
e2xTV3Y88DrVk12eUrsvMgOK7EUAYO0fEKFfNvWA93qjzm6I5qJzx32nDHSTY7Wj
CSvYS87q0KlHho8fPPwZXTWy/687eVs+/i8n10G+qR6cJ8fJo++YRW4KzeGMIzd4
TFVRW1+FSVFYF5O0ckIA7UMJKfSkGpdVM5CaJiJR4pCvjCdnWudvqgguaR2QSEr3
B4ur3eRWYq4tTLY5I1QoXNB4orNV5SReuyqqCyzTuho8qAmw6EMG3E/pr670fs8M
YEAo5SL0uOCnefOk0LyBNNOsyK05XPSoVNQ2SvMekPpllOO/Yg2AC4LD/JEAr2ZK
ZqWOeoK5dKB2MZA8t8oi4/fKioQTwon6o2NVYRjxgOaFi1vU96rLoGDq2Qf5WNkz
0FT4gZzdNKGA/C9YtOju/zh0/PWbqwoY1418dlyMOQCM/S7dsWERUl6UO9zDCgBi
3r+6A0Wpn6y7mFNLnBK94MiulHOo1/pf1B3yy72DVDx48XfwleahNv5O3bf/XWo5
Qp11Z1sK1RmQvZ2LAXP1jC4bf23D3OPL85gSpv6PRALrXBkyjZYRwcWYGH4wN/gH
9K0As4P8TtbyvkdBKCOYeYxuZLRp7+1mQbYaE1YBAT5cz4idI2vTc6RIwD39bAbB
u9t3V6O8YCqrCyX+WAoXWNd/l9LTagzqdkjXjs9zkOLcxmveVTIMNREf2edvPB4V
IRg4+Yi+UC69NJyj/2RFrLlGUPJ4yeNI2dn5DNKznyI/zHbfiDNIDexkvtDyacYi
1cqgo+0zFjH9BHQvRMtnPf81qmQClzP43ZyddhYqMc+w/MjEQZLqH25G9TAsk8zo
XIxQ6GD6PUxgOoFxYHwITN5qH9xFju5YtuxjCg8t4Tz0iFsUkbucKMFgILgNxno2
S0ZZYx3jlcY9g+dVbg0Mmkedn03QvoId/t0RiEwkAluiESaHF3U3omrJ2hxn/zAA
AQkB8VWS6JuutdziXpDTn5QrfgwYqYEAahjHPUUTYGyrQpryN8OHCgE6U8BxZDSt
c6Pr6rTDSiWDwh0kGzoe08J3ObKQ8jS7c/Rx1wiCLNYVmPik+rphvuEWuTSN4T1H
BUp1J7olv9yTIh7ie1Mk/FgnegU+irDlozitFv6J4Z/DDl+dRNHskpFQNjshGNJy
WjNodlmLUggC5x2sJF5tpAFtX4KkvbFUFT6s7JW1ZNGt6Ky5+a7/BnbjJBQQ9YnR
GQeTSJ2gCLnybVlUY2tmc/mh/1aUlXR/QXkT8NWc/r0k2BKIhq3ELbKBu5p3hBcy
4FKnbvQIYNRPMEtZ4NX6ZJWj9r/nvpcBQijpFg4aJTzqG97ENn6vC98DhlHZg/nA
IBzanHj7yXfeIjcr8UAlTSwoNjIsQh7sIMhKygf0MPusU0wxQyighJWWUY2ioBwS
mavdX10MtjMG3CZeYESjOkGzsG36/xp4WLhG+kJhmgMgd0Ei43RNInLb7eHgBBGc
RtaFTPtC1PEYtfcqs+fCINrkajH4lTvylnty1t6r6T2pU3rjNieteDXZCeQj26wh
WTLvBSDBVOK8EMWh9LOpvpUo48PW/cUqolZhpYGohVp4IV7FevhnjEdFYvdNy+ix
cOPMTIKxuT4CwwQh2B1G9TmZxSptQFhm39fdj/4rGyP0XbE2V+cuq7aYembwTXWs
FszKGF+2TOlKA//cDDIQ5IWzSb1S+lqbPRJzF1AJpzfKi8O62L1R3WP6XFj+BWyn
M+htd+TLxmw243JgFT+4YzCnN+uPRhlO0iTqroBeSgfpF3vbRcOYaoG79jLv+BId
Zy+UkA/GYhJiGalYI7OwunaiOYdj9JfL0tmrTybmp11SzyPjfP4UGsSgypE1wYIU
Tm1tJwEY/zUStYX4N2lUTuFMsFcxSzfh+Yx7DNRGN+neKPT4P5mBf9aI+/IuqvYI
wUQ15pwNVFNizF7JpDv+L22KegRI7N1AqtHpQbQtd8ijMsDpuEHNDJJGwkdozoEN
tLLU7jQ2KyY35wewRq2tY6bPjxJegOHpQ3kiANqIEZoclAWGnGf3RXjP9FbNtrzI
BjB/E7TmJ6PQCju1+/7cwpvBFYFisCKKN9qvjtHpn1tY/l/XIBIPNHTIPG5jJQ6c
hRNdmYHoLPjnVfcJ+xEGN3f9dyyjuuDcXRcn1hOuPRbQren7FkKKKdqhzKXiFmm1
1Ajmdv/nvCHsS3zAU6b1LGmqvzeQvlZbmMJje1j3sXnSJZfkMTIjfSpqNbNKLt+l
NAJfpKJ/peZRXEo9p3CjOFxJoCKc/IaHopF1TQF+AbqoU9fG0g4bzEn5TwFvjcCN
+yQ1MmtDjHp9uCAmQTpoATXEbQ2mxCmI6lwyoKJDP7oVkHdX1hGKTBh9EYVI7ZTi
AkfpJfiLzjipBQ46/nhmZiMfprYuIWiUrp6syk5d306Eli4VXbvGtmyY9vf5Q7LX
N0MQ24SA55/1F7zk6IdCVBDPHMuhOLeF0vc0LBJa5I/UYzjstItCjvpNl/efeQ/s
ZgI+qNj77/6kVK3UfdYzdgPA0hIjrhpZJ4x6/E/OO4Tl91CZw9DSBAoKNB8m2Ljm
+ejnlmmi4MVLHIJ/67El4ZR5ZlVDFPxuS4BT9CIuanwyy+824WYeyAviIJjumWCM
JTuL+KWO9lB8G/Q2aEbGz7DKWe/I6fSu8SASCJ5c8b5gZ7q0GX+0k8vCgY0p2Zd5
fKfwlGLcg/6lxot7t5JAVOZmPXXyyV0GwpwrZwnEIensmSR3HTaqwvDm1gJTLKti
q44VoWirKHPV6MncqEKWjjJwp9GZP8bptwhV/OazIEKQ4Nidu1TeU9l6nS/brtiL
Jj1I8RMvh8pmA/4VSSEwqmfkC1fs62psqHakYirh911UoGQKYNq/e0n7mEctOGht
le/ZwUP1Ka3rvnXKuVLNoBDnmaCFyElRDO/R4KDtZOENbuwGMukgIrlg+vPD/Fz2
yrqgENlU7+8GvISdtSZyUhcNfnzcVU4bSmKQoRRlyaFsUXMBbM/gcE9ZLmLuyU2W
KOyUclY/CR7JXdkzYZkscZmB8WzXKuC691mCY2U3NtPES4SZamvWbuRYyzHwL/qQ
YOtz5XWUEn+3kVghFK8c1uleTRZaDpHY8G/zgAZmH70PFfL2wqnsEAoOtpI9jc1X
8oFgx47d+d9cLoSuOnAjGaIGTJ9quUVNoYiwagmVoQpRZjyeb8kyptD+Uz5nDihY
yEkyYbN6RE0PRiedymrRieH2UgGwB/ah86kokkH9Z2V0h3ucDG/6XK5YFdxr8nJA
vSm59pDsK2vnH80PpDIyHguNPRvSFiuJjEGOazVFj4RyJ8iRmw7QyKrr8B4NUf+M
9jk1mFmtXhN96VqcDTAxdGNvBl1ly47GQ0K34KlmxnzWygMltBXwSdREaSp1OnYS
DjMIHfzp3yMf24JGDBex6lzQkVCdoxQnOFByEOHobciAOTiwysP1U1mHE/hF7nNC
Vmc0q1lV8l/xvTbw9r5kduY615I3ts+JWZ/JvuSryYfr/KTkl9Uc/Zm5D+wlHa5V
jyyW/0XCBaxe0Jyjgfz4pP6S417Nfjw8intpQIfEo/lkrWzeEyJM/Mhw/hP7R9bB
T2an5PD6Grxl3xo8Yp8Mxm1LPXkV3lsUlLcb3+dEslAD4tAqs/COfq4jLsDyr91D
dPdCWnYkAXOdriL02XOOK8ifTCgFZEgrWGvGVOlOUs7hscOk+Ci/h78HUILnBIAh
7ERYsdX+6yWZ30HiH/sIerFiKVR23/8KRw88MEFDctyyb5eCwZIz48mzMupHQ1Vq
cjBeUOJi6bBkThWsw7oOZyBHQrt0U524okJUVQjdHtakwUkmXi0vQKkFYENMGbls
D0kQ54frfPff8VTxTLacTrDX4uJSpD9risv3eSnY0GSbdbMf1mCCb/3C3Lboyx6O
EXKBN6h4wLZ5WGyyRqgWpvba5MacbWdi8tXO1Vah2DgwuiOoQ/DTxFXpucDCHsK3
Pn379RqssXVMOo9mrwpoEPUBbwiBvGljW6qaJnVuwdQRu3Eu22Pl2CRaYUR7sImR
chmJczjRrfkgI+YCkLCHAC1h1dbc6KPkuzjTTTKSi9++Npq4bg7H/BJibZkaMSDV
FsCSlFW37vWwW6WCa4WEhybRRk4/nXxh+JVsEGAtKhigm4sHpCHPThSFcWbCKMWe
dw4qCPyCjihHPOlFnxIdU4fkc6ksozDvjRtxyIk6aFwVjmfLM+SDOjT0OIYzS2nO
fsOFIfysSVfHotUYN0R1QPvhMVqOwlRXHaQ00hFw+/hb44v7/MKloN6c8e5q0l+A
3eUo7AyBmPsyVcs0yynJfTXj6VkBZnVJFqvQBSH5kC+dPvbdBf0T7Sfm5HutHWqN
v8U/LXU9WbKx/9QugMsVF2O/vplw+tNLJFHBzc1meSB55zh+nIpntq7clEYevd1W
ALGyP7WaIhAuooINL1Q2IrvHutDCriHHPUFxcP2TZ4UtExg3yOOS2/sQiAlkBo9o
UtNJQTZ8+qMUW/9YDb2iIo9CLrIVmicZ+hQRwa4FhpNsX1xk99fzF/MI9s+nqKOS
DGog1kBEuqxEIrXT9OTs4l78uh3QN8X8cWCCFRCuLUClg0J+rWTzGtlLEsI1Kwd5
N7e1X6CL8onsGMHHQizgDA6EVZhEzZSNK/GHu4J1Lb2rX5pOAnLbY+OkmNO5x+mV
m0p3japtta0F9a4YqfLL3DBqwZNiCcW3FT+YNOPdxoqHTF85yw7skdRPR73BYD1O
xrDq5bOyEUkuLSQVAuzanJxfkujCPfU4laL7oOw08NIGCmtuwA13JKg5UsogT6cH
2PXNA2Jhyt1mOqGZb19+QxKKa+RcMYKxg8EwKi1dGdjnWG/Qxka72OiRi3CwwPdr
8U1nPT2TIpWO/mBBiNpkpvP0RM0U5hYWAD3Dq5uJOfdpIB+ucRnqkQtqf++fdElC
jr6xibh8QX92rrjONukKRQCB4gcuAb/B6GeDFT+v2dwD9OVmsTz1zaBE4jNmr1dS
PPWGZmezNSBUHUDnMaJo7Pdx5aP2lxeCw24ZxO1UE5JT0g+Q6T80/WWklH5OerHh
MvmF+J2JEmH9K3aeO9MWsBpJQWWzywp6VDe8QQWNBDVymMkByg+UqHRiIDB+7+Ib
f5gunumgVXAM8pajxvd0aechQonWngbegRvu+gRIDqM57gePEHsI6wHygRzVI+Ip
eFIId6kZZlcel685n6q9FOS6aRIK43+lyPDsRLZ9IDwGfRkNGEtWPmokOSj9Kzhl
2PMAu83JvCUJmQxMAq9HnKujwlQgJkLXWm8IoADr+8f6OiTEO+pCiyW5a+mmQsJ9
W8qu9KaEkQPNY0JU66rYbEkeyHFi21GqlfPZnTsmoBTzIjQQf8oGjCVOZwmNZ54I
oRC7JGFzCp6sNmBvVb6pu8V3nGooe2+0DG590BpUSoqW4N6q/mNpHCWFU+nI6n0R
rHAddd0tO7o2uXeTj4yTZs1KMycOtbTd5/S96JL2TGOnfSY3JulTbDDdd14G350H
b6OzO9uPeMigrwrrjKru3WqeXFri2CAe/moD3euar7x+wCA6wpgEjctX+faRJhEn
C87a4U5pqmtqfYVxoynEx0K28cwIw+jVWEc0ufUW/UcYoyGn+X/pgIf7Fyp2eHy6
7j28R7p6EKpEeKBBsiZQcOKYDmPCaDjbmgqkAnFwXWRFMFEhTmFhB165Kk+H/Z6i
0wMDGChqCCr5cuaqXvLh8tssPomIAw8ruGkDRv2sa3L3fwldYNjc35/qYKpPw/zd
cc2qnOgjtwFgIhJhUns3mByJ/L3ry+hUDOCN+U9cZC9EIJyU2IS84yllKw1wdHcX
eRjhV60l2N+kVjLMtH7ASScb0bm54N8gLyzR8H1nvxdDnS25rhx/XQwfWpl6ZFnm
nPKO0EUi5VAKRAFsgFd+hESiiUYlU44BkjyJo1GT3VUk+ui0VLRuo6YH5CUead7u
8m/AIfGkyGMFNFIL3tu5wdy7iFW8wTaj7WWyQReuTUPRjvyVZwLF7Mncjkzc8Gft
VooDjAYnyH+K/SRHNnC24JsMtD01/sfWKmTjIH3cmukrHRj4j7Ozz0WSmdge4rQe
fLgOTg8DUni2V/T/8b0+Pzv8amztVCPgdy/2MveS6Ctk/OsdrSumHEtlKxu5n/5H
KnBLwu2CoHzzNc5J8oRUR4PCQxGZOE5SgXUOjViSXKyP3ywMmSU5m0bbDeRqk5gJ
T9wAoheLrdKEShbJcf6JiAJULskuzWDKN7Jpab7OUbA0jlmXMcwlFveF8oJS8015
vP2WxaD+PI4jdZNZITGCX/1AIsjUGGHL405bIS5k+DTaS5/OLgLqB3euZZYmX4BL
jKR36KTngfqgggw99U97bg1ths9w2t/i8bTSGxniN+VDWwJUEpNV0Ko7C4F2yRGc
NAGIL1tdfBrBmLg7PjDd9PQftL59knCxlSO9TN3GaeWY/6medPVYxdYL9xtqDJ6U
Q7ekTd84ST5uDyARh0aF5/2fLp/WIpPkd14imwtQaJoQaqUuEDem1D/zO1HHMm4U
fF9hdPj/VdphY66ks8Q4ijQ4jRMEtOXOoQ/X/hHTBo9KaqKdu5t247csY7EQ2Y7A
WnoQwtd4/yohpVg/kcvnxb0TDaFB5yxLVPu2rI9bufNcYyW3z2Q5nxnRsSm6hChm
X2BvTFbd5/CYiaFRGP1t42mWcPRvdeTvQChnXJDKINwSTCpDW4dg1TOklA41xYOX
/0kudQqPMp0IiFYjykdU8/2yInPe2m7zIWhJUrbM/biqQzesUlqWibRb97Miyycp
Ch1QK2M7gkvJHyKTYfLB6jiNNlK5NVf2AZ84Z6GEFRSf8tTNkWETTjhqhmuXao47
MRQcB47Ew0iJbWv0GP1FbWLe8mf/++wnNK7gLKScX6F9rDaK87owMOlvyvgNL8kT
efVlcnd/QlFMt3R0qPtoJtvAuYG4XQ2BJXtVQSx+68Nawtbu13acaTCCfl8n2zcB
YsK+LCQp2J//8Kobauq0EGxp9H6+rzGB+7S1xfoFqmTkYQhBD76wx9Nfj7aPvYZu
Y9/d4+Aq0nw+zGDdRZ9/J9IRcDQlSlW1XTsFrlEqsV9laQZ949gB1G/mpDuH8Fdw
H/RozDmGDOKyyKFu1BMoQ5gCnm3K9ros3zLIokiOKd93SKqSqJyR6W2p9ja0eRr0
lh1ACHlH4RNEQB2NfxGj/NsMjRCPtsFsq75dfGa9AklCFSWL25iMthk/ryHXEJ64
1d0dLwcXLfIz75ZTgn+uR25broL857iXDGAffwiyuRnP3R8bg3o0CPHRUBMKvVR5
JL/yxx6zlB2tsjyiGWcM5LyRN+w7Ilj2aMjJwIQq/UeHsuoA8rs4XTT0qLebKKsK
YZRuzmQZfvkvZvewopKksNbD0XOMVKNBRfo8KGW2TWPDSN0fHjG/o7wsuF0eQmg5
2S//1iGw/qQB1dRJ5Uq++Pt0u6xHFDX2HCL6eyA3rNf/jGGE94gm1DXwzqt8iSpa
5pVWXJlMPctxkwOHrycNmwMMpr4pr404OUJgz1XIKEs35JNFwJ4aMYKSH60Lf6HG
lDEKI67dS9ZTmyTnLvbPOqkpBhfTm1gX68HOh9B+3q5u8OLi/3C8QmeNbgIqAgrw
r6OVHe/5vxOXYtudF0/KlFZQkJC9R9UVHspZ3OHCSHyyUlIDO5p5WrNicuS+iPOO
b9f1Xjp2AtI7rJkIKYYd/evCoFDx1W/FmBfTrcWMeivonmcGLBQAb65qTwu3i28E
ymsSpSy68x8MzM06osEHQqVDYFfLYCC1Gi1TBzf/OeDDFtZEgYst2G2GOnbmLK07
Eb+an2PdJlWTT01nT8DJqmsu6Cz62Kg9E0XjM5UtsoLKewzD7Usrb+pMKlIUmCuF
PnsKcgFzSo/hidKdMr7Mh/w1sAhrP5r+CFzHjs0AgBKQhkGlpTHtM8niHIyuZbtv
7TOo//Mh4H/67pwQ4rqd8IJjXuuMrpV1vm12wx8947R+oyq8l1h8tY+G0XWVJ/Y1
6rJUEFcWii/waBIQie0ObFshLuBlrK8ResHaKkS2Elznfie4uae87nl8OpsZEruU
HGf0jjuP6yHUr0xmvNS03DfovClYLqDqQEhxEliUbHIPUgwUviWZRvZFi/F0Lvw9
rTKtV62KsB7xDLWoKHiNhU7MX6V5PzoKRq7FT1etU1z/4oBiq+g/f9v93Sj/3qmM
cNp+O+EngbmJH+lKamy/Kywkftn/NU3XIiU1o8PkEDmhbD9bWHP6gBS2aFT27v1V
A8piRn/pv+DkW1h1rgFKnsMIm3Rhd8hYc0+QfsrvmikNZW281SpioaeTZFB66IQs
8fDzckBu4xzjnAUI6rWAVxuKhRNiH2QRKzHzKGe2UcVhlArt1rvwDsNiUbg7CyzC
9/+D1JYMTvVpg3aBYeNcs0Y9BSPnt+78+b0Mel8ojHncLkDrxrJ/3KnDCn6jwkOv
qqSOnvoq/STfqveCdJSFB9WDglGMvcWC4bALvx5k5KA7+zkIv0trli3lE6OvZRYd
YUfU2VkUQ33yK1wTLJGkrSNZypbx+0xP0F4W1X7ZwYR/OKxzn17K6S6PxnxnANHE
27JZHoS8NVcmuHnBx7jBodLAw+7CHdSPxaK8yO1JJ/Vx+RWCpyH43La/O5pF5Gmm
byvTQPs4I/Xc5VqJt7vi9PK5b/A39CGUH/oA6SJitEY6iI7lqAmXHh1tszkrkO0J
FFy+Elu04mpaffvORF0dOWt7kIZB5uDK9zE79DisGjITmdy8A6eJZaAXnk39dCY/
+YKema0QEMw8MsNjNvoVXD/P+eh/nAJXJFPmlkyfXL3bFCqx047gJh0OS/FyUAim
n4co+uwsKwlN8IQDcVbXm8cXZEXHMPCOKphZGyNL9OAm//S+TkK0wjnZJNWYEdmE
U+hvlj1uasMV03Uv1zEuDA9AYEW/ZxKH+lI9LmpIucNZhMn4XAOR3zAw/nFnPCSj
6pmZyKiVeU99xUfoyqtP4tvMmbM0BpL10z7KjS+yGvOZkCOx+eSh3GkWMSJ5LIyt
oaUAbDbo+YCh/uV302zSNWkpWKYDrYYSbxgTQaf7+zTprfRJh9gwnlZsKY9nNc1e
ohDVq7jBI1kWl88kg51n2tQ0/196LSKZRK+0AOKIiotk1bBTYrTTpeK8yl7O197m
03jZywS88Oc+H8U4+042jOlM2l8fw2d1oRV9pqeDvpBfC7NBgJlT0f0E49iQc7Nz
2+sVcnEGbQA/yadNqne6d3RY+EVF8SFS3Wx3J2aAjyOuoZWrAGMrpQH4pPwNkNeX
rHohUs02bjM3x6lO86JS5I68zJ85O56VhP3IQI4NBswbXqDGZhzfxlYbht3JdDQy
csF/es0KRFSKQkj+UhSUOHEqLiN3YLJvGgNqKWpPxG2l42WAynVUXY596DBjz7vF
wOyeW6rUDntqE3JFUkMQHm3SZhF5WAxpchcaNrW8zY6J51F+RH23ea6f/0yrTyDQ
vT92oXh4859SgZlINBNwiIvvxkTUUfUimTI0+RmjZTxhFh7FViBfl2hqojYfq24o
6D+swF/lQEAcoKUZMCUsjVuPp5P9OxyArM481478o4i5YyrdR76wD7lxizNWXbG+
bAq03eNxv1bFQUFc292NIATVcxvzv1kgIqRCNzaIGhkPxpT8yH61c0IN+K9ssdHQ
5XDeRX5Q3Ywg/+oxoc7A7/roHhSdeh3Umrz8IOjpcl9hawDsUw6LNL1RWIm2A43t
b3uN93Ao9KEE8zb5ybt5GwP2XzQucfQaEGNxURpjFyYT7ZASeJliOisDywmPGjlH
JR2JkHtlLhehB/BdpUUQEIJdn5Q3chElztOVSLuXTFFVxQlzeakvlLDU/NoV6B/B
p+2jV8dOOfYRCdd21zPuq1GR/yn0f8030OWhF8k8WOmqCGUtFrNW0aqs3iVaiw5L
p3BTQFn3UBUbTWL1BM7xDZ08A7pr9XvaJmEshoQo31GoTA7HhwQ8tszePluwzuSh
G6+5t5rIq3NuEN+uiA29oLqKZ8KKqC4e4Ji/c5pn2QSybD9qqVMae/n71Y+g5T1u
0PWoZlkzO1zDwDTwctqeGAFxVK+NRWkEtNHu1HACXpVYh/BlJMV3Xlw6Z8+I81r3
tqPXrL6recLskzj0WvgY3KykOrrg9zG785CFPRgv7o3lcpL1SrbSn+h1trVPBVDW
VCDgrT6Za0Ibi89ikFMU9hhouzE0aFAg2Z9H2W9ww8URvhNIWsps5j8AMczcEZc9
WSCTINYD0smmN4mmsJPhEQUnsy/HUHunZWnG++diQdbx+zz8CY5IRuVGMdUQ/4DT
JEikdIUOXFfXXTmBc4zo6We9vwcap8bnDdqBqNHBNo/4xgiyzDZ7Ea7wo3EiUXDG
txrmw00tpQ1JE42l6j+XAT35XfmfEnDI86ZX7BKMuY3tnuwEohSNjf5W2e59Q3pj
k3SFBURovZpbHpELn/Hr5PLQ5Ap8m7ajjg9TSuL68v/Nd9sGzi2UJGcoQ4GxexQK
i5KJ/xy/B91rfIaIAm2GRXQhgWDBoGpPfq1a0cT5QqHwxUEedq/dney/uEE27B+o
glKlZkeYBTZFdGT083fz9mRmwgpzCVId0IrKcW+iR2vCfR1Yq4v6PDhQfFtp4fSG
purXCPDP4ssPpMvq05O6bv+lTIe7+WDbXNZU9eJXklZDGThg+hTlAaDlLhEBpcnO
SNmKPkyI08Dx622/Kv1FS9zj6HvdW5bnqs6xvktdjyOblEV1CsRNWe2ho4eAXBBn
i9lDf8+BAXGkfH8UWS9yzxosClvFU7pd/Y2xn6nDRsnQhjVnBT/hqzfbXAkbMVx6
A1kLPm8oRbUdisV4dxiq04tks9TxRAmQTjlHgS0vqS8Wk8bNy45Rix3tJkAoz7S/
FyNGnNqqKjWrxB37xusPnkguk1fxFVK4hcwSySMuiYSTED/hkVmljajqx+jeIu7T
j3CXsA5OcppKaTnT08nnZlcYzcCNFfuue7BBS4u3/THtctTItnNS9LXBQEuZHSGd
RQAzpPPPn3Y/KEG/z/i3T4C8QT2aUaPikNmRg9NcnVsyKQuNHqWACuc2ByldLtOj
A75OZdT0puFztDZcCq5vJoCixQFVJ37hDPi9hA6f1RIrtJ+jtntenmtFU7ypAcgc
FvFrFXCfy83xuMlLGLootGTmrzZg8h/9+nKa6dRyd+gcCt7OeB/rOJWdRAyN6UU1
DUdSadWlg7hPnjHvJeCg2mxtxkGd+oo5BUfu5q9x+Jr3OwSMtaKwEWgfChnWEaU6
pBDVxcMCDmx719Rqq/ndjQyJpWXBGZ0N+iSOlPNToiPAD+DZqpj0cOg8bcllBM/L
IIiOYr15JZNcCO7eTY87SO2WM1rH8nZURLpfFPry0qTo9lV0z9zYoY1WVWL6IkoJ
8E6u8RHNUukmhOy/eHb7c9zb1OTcM2iIPIcyEXqhd7MQ5owtYmkaHpAB4IK/mxbj
tZFFhToPXIPuKleftes8Bpu/jhQ8cn/1ftjgGWmC/3B2Rq1M3sCpE56Fxbu0eY4+
Cq2xqr0mPjPDU9BumrTb1wBavUuWHoo6UZw65aeDb6FghU/xg+nQiDL9UjK0Lba/
J/h0pCchI/KExhY/Cijw9dp8j7Jk/Ppng+5SYmESg0rWDv/mtmoMfLN9/Gz+LvIO
wXuPm4ylPG4vHkNdcCUqu2Mk9PGdUNVquhx+QmXAZshjREZdSd+MnlDhTEZJIGFB
Eie+ckUk7nP67NWtzwFwdUA4dnhqHxMhcB+ddw96GFEZVSFFg9bJRWk5Ru2IeO56
vBd08OHpGx9DjiimZCWZ+BbYId2kfU28gVLDZhpfAQkul1kraQFhAcoWdZacVLAH
nIjjJuZzv/hMAtgtY88RH7LCPu+gSJo5vamaQ8XbcEQWsSJI1QouFMKFumlO90xy
XUf9bprMcBQ5v227paF8pPdwoFiIm+Sf4PqRyTcIyNRB74WWmI8XRVMXiy7rFKV8
RDMpb4o6f57DJkPWeSSkVI/OZehhbJScoEydS47xnUE15aE96LjbMOm30oTSO/hH
0levvQLL4sQvNDPxM00emv6mIpyOndRkbcKNbBFIt7jALZnCIWATznrK/YkPRMSe
OjbcEtItcN3hWwivqrsBVKfrqdBHTDyFLnwh9/CVe3IRlrrAveJprA9LepkZ4H+I
8mHi0HedCIext6aFFoRNELJy6Od1zlLX5xutheN5l1/6Z3LsW2r9Di45qKDNiAF5
/NSqVpjq9ePL8RkA8KUUyODjXaUZKSDeGYawtkWWfW61ab4TqF46TSbfnZ9lmxvI
Jm3LyDPIZ5DVg0+s4jbS6DfNGMg7u1DzjyYOksnKtJ7Oh1meBtf0oFEkX5nOPom6
saebylqV+r2/aXJRX4duh45v0F/YsD+XHVfOufy5qiv2qaa61y9eRWPVePq3qpui
+ik9rNw/xYowzorCvrKXdxEpQUMMcj5vN53JHTBFMk+jj7dh08HthKv1cp7jS5Rt
KUHIMukOuXsQjD61ho0flWYCn3ZfxgogT/gbuYnGTUG/xpE26IPwHCiOeZ5uTNn9
oIeG0s93OeqoClgg7ZWOgV9aGNRKpGlY8+y5oA6wbSYyGLdNwGfoukqLgr1Owv7o
hc96PHllg3h3V6lxmCIQfkWngH0XHr6BOzeRws+SB+u4+mXvzZVgAAKTAHQHL1UN
ebffDfV1vLtCZC7qR6rf/dn0u++mP7WrceNE/ur/Q/9AzP0P64UcRGfs+IhuLh61
DRvb7v/hVXlPedzTwUF+EF6MIzw9V0P/Fuo9IA+ilbs17iCkugjeV7Azv3418jJY
VlBDDC+4IO1i1IcPCJeile4xzQ8q3UyGx9dL76Q6fBLCa0p+gH1U4gdpbVfzkxU9
+WYs+qDw9iBwAcbnATLUv2qPb+CBDJUZZjAIRAlJSWTWlTIdv6Ys6EqM86AlV9Qh
/TLiihXM2Q+nJC6Hka7mOEXb/1uqcRGpfvlOLJKx2j30N9focBANKsrmmPo+Ovno
PWTIhi8rZEfbsYIAtaTveUlPH+ZDb55mosS63t7GUp9U7SezUrrls09FUUDgXCla
ErxJPuVu4nGDjZnKALs4Q6P2y3V0tlFx02clnhHpeBDE3gihoc1malQ3mdMbA2Gm
XJUrlrMMhzlil3o6Ej7AfYlsfE6pYgg6eTf1QNBQ1tnrN4aUK+/gRH4M3GXdw/BH
3+jq7oPAmR8iZtCz3KQwpnfsgjaLv1ffKb4qV9g3Fc/Zd8S2GheNjdEh0GOTa6m5
ev8a1Rwb8kQnmk5xtbMuQN8xYMiaehI5wIrPmKuCla3qSbIFJEVhkzT0oEUOwH6a
0g2g3Y6af/RnjdFf3x4moI+/xGhVY2LpQ8HgikZmoqH09jVF/Uc6QRppxb1PXDpy
AXPIXA6XJlKteW441u/QL4cGDR4KYERCKSi/WdZNTI/iCln0Y4AAMrPPtp/G32r/
RRsjSKmSPvzMnsZsRjKvMpDcbJ8yk84uh5SPBaC0CrTBFAMZ0/Bh18quc8UqCpwH
yFeeCw0I/PncxnTYoPGLoyZeDec0LxqHpmdTOD8of9zGUveQ3WmiAtB0dDyqAdVK
WAZcXIaWnoQ7cA3RPR4Ui5EnqwMteEpxbpYBYBgzZrhexhqa6Jmf61juKCIRKxjf
K9sEjXAkqFf8sRKCgJsr5LTCboZomC0IRpHco3uhZr0M5lhPdaTnoJWzar6PAzdh
/CUkJzVqUrlKeJJp+VUq6/u8+GwuHjgO71bD2nzzA0DrsqXXZS6i0EueTTvEY9L5
1uFfBx9giLkapRozPxcdJgrY4Q26STGo4KQ68m3y6C02FwD3wE6cZQoNqquu2ew3
V7WJiqRw5SCZlYD0hr3jduU+70TMqTzu9uSy2zjKGknGgg9HYI8DUUdf4hZa+ZUQ
t2/d0971OaJKjWFC5PdCwiAd1tUTx5l6gOcwVOeDnLXxiJvCF7EuTnwa3nVjI7+i
ehtiF/xW93l1weovZwlV2BXeXgmVo41WT+RjdGGc25Oysdt7WJ6fih3TzUX3nqZL
ZzZhMvyr8HwB5qi2qQpG4E39oUwz3dxXLc0lJFN+LOiPQxWThyVYVbyMC9sdgm9W
tzTvLiqNvze6VmithGq1NoTkzOfAABJ42rWRjIHheJ9YgHPgIgpxg4TuUFtqHYbV
d88sZoMmkgBFRgN1g6PNYHxGX0JFUpzJUEpRxjmukIo1qwTi3Rslwa8wXDlEKnco
/pDYga8aWIdy0tVFG15MfcLbhjDorikyoAtyQgXZhVWGdknInsNKNp0mJpJfru7H
E6fWYj3bXhZKq0WY5USfQlEG4RetDSwg5nQrKEJs26KYfkan2RI2R+igVJm/Jdb/
bIF3ADBC6YI/U/dI9Y7yPw67GuuMxrChpu9lS+4R4e6a3O4SCXv92rqsRwnLUfIv
es5RPYXS0SbNnFRDXGc6gl4CtIOFDJ/jaFQrY6QhfvaQ93oUCmWI1boWePMlYyDC
gr1ERT5AFEw7AKl6rOZIhDjBvGRA9cAWUUnMN45dCw1NPRBXexAuXLoCwIaRyFs+
M62nhVlK8KYSIkdynkYlYxObtsThm5D3LyaWPX4f/QPsTXDUkN6btEsy0MXI2n3i
B+loIfO2PcYgsH0ZETbp6ma0U0qyh2j9bM2afct3CE3nRsdFarnurot95BjemPv7
htmhGeb1tkjxPfnOANUjBPA2LYWYsHRhq1RHLvhOBs2ykKZR/Jl/AZR1KwLO0J/w
T+JKV7Q4uBBSjjY2q1IH9mhj2hZlQQ7PkesmCHAUy7fRJ+/IeDneacxbVL428/1v
JoDnml+XO1CFwb1Ja4wA3dLqcKRgNwYO3Y4v4ddNQxRI1REXiSuWvOCfrcpVs8qV
S2GL6U1MZaJd38wt8h9efErZ28KLdZc1/9fa3QI4mOUyrYpsJ93R4S0OhrMUq9XY
NYOk9vLdfuUqeNnMcnRQyXEM4iLYfohkgZFhWJUpZ3Vwc47F8VoRKMx6myZq0pmL
hv916r3zJ38f9SmSyHRF1/sqlge2dK/oXF3UE9vz3608PaxHwgzSJQWUW1xelRER
dKarHw/3ynJVEtA+U8j0UekhzBuXrrLhcRzAN9KUh5YFTs3TQ8AD/9ajnsKft53A
Pu23RExPW8jHYkiCs99UZFqsVRgLm8b7gn2koogQEByfAfXGSBv6Fds1mLRKNvBt
sWOOT0vhnngXvvko8Sd40MxfehS4f5s80DpgOaMnoXODdWhfakthTrmG0hNhnBm6
snc4gNaFlo+StQAxeOm4Hx3dQ71A2xIfGvDMLm84HVNbw1Ojxw//a9Qg4ByAdTr3
yW/QW5wTL80cioVEcjWd6WPYxYLe9665g0pfSwMoJfQC+bpqqmbGmdLpl2G0FcsK
3S0/+oOO3hectFvOYpaw+rzr/Skw8A5o7Lb8gIuiDkED9ihkQS6GMT+QsPFggvPb
BqePTzlzYPbDKTybV2fH0pWT7IL1Vkh7RuItE0zlXp/X/Qax1OhAOnmCehaQYynw
/gVaYURVx6d3rMkyA0mT/DSDu/P86b4F6cYTjU15jvMOhc9X+DJZd0tHoYlCuxdU
SnakdGWbQkfRJGCXYlff+DUhMeLjVsOw0h7O+omFTqB1MFbM/5L1mWTHSYJrKQn7
+9FknD08fkBdAWMdKCuLi8Myu7EdJNtAFQx4plKl36wtghLz89XhdL4euZq5OWwu
s/JQOcBD5Hq4Vel7Rwkx30D7euQ1r8L25N3QBFMidRWL6j217M2GnDJRzTyy4T0G
eLqKdUhNQ/EQq1SgzMgB3QigsMMxSK31WQ24Zds7VBvdFOHPb0MWX6QODoDGEl8F
0bpFlfToZ5O9Vw2HgLq9SqCbR7t5gw2kn3Qsdak64wzNNdOrekzy2D7p8VoDOO4z
QcYRDLxgBYWb8t6+/GYx5SMh1Ci8347DtXJa0sEVAuj4y/EXQmxkk8NOMeOfQeWK
4mQdF6dkU3b1t6K1+4bI+Eztq2gUnqwFRhcvnILbOGIAcyAZmwyRDbCtOlcwPlV3
yGM43ysEWFCYGGICH1N16OLzKkX1IVK0Dzfe4sQSutaAGFqsM+ap8lHkauX5xZwC
r6p8lbsNJvP+bU4WLfAM62qyiE+dCEJNqQVOxZLs2ApFP/X0o4Xs47W7sIXCERez
dl99KjvoX4N5lkP8g08Jwz1TkK4KjcWs5IqBWmxzS8+q/bRac9ErO17a3KTlSQgS
wpxfOFEzV6MxaDs3tXJVrF1IUuA7dNcIwuXcoXpPeu1pNiT75yyY1Dbe9bDx5wMr
WnNdXv+lQEiy/IdnwfNQF32ixCoLjzI1NpGQQGxk0VVdZe4a1hhmP2W+KMIxN6hW
6whlX0oPVN55QYJM4/b1RZiew2CsAbWS0OXNr5Qo2QxQ0q0yc4A9EyxSKbCtzO2g
thNk2mHAak8HtGN9RTphNuoM5d99olb7bFiYIvuaKa3nIZcLmwvi2OtXp4ELMod2
rEMV4w3sWLwP2etU+b3qqzx2mzkpfvyLCR6eZB+unMkK9KSCDCvl9pNA6OCAvOAt
Kyii9/mhE6WeyTaAOLW387HeAF7PcWwAJ08dPHFBAW8IG4tQIW+qfIywDXXasICG
6Rn9IvkGKoAETCfVq68oxa2MWkdWBwxjuB9gRPMBpXIQtySf4LSsvjjGYoVOO9um
B5WIFFDGxO3M6FlupAESeTvJ/OUvgjzLUcz+StrmywUPueHoaVT/SsCqFNGTXpIr
ISh3aRZQJLN7ueOhbXnhEXQElImEaKpIPR3Ch8uYxWb6JgdVaeqzUMRwuxCLlmo+
FBV9UuFntdKW2P/hq5eflBMDK8AH1+TyvOuZ7xB7inWaWr6/kLj5HEThjhBf1e6E
oNU0CD7gtoz4NfT9udu8/J77MhMj1H0qolQzsff//rm1l7BfibDd9a5lAbeTHwep
g1L3Kg8D5Rn9N/hvwyXpMPMPeEV3KQyCAvSoz/7e9DpwHn5pIY96p5j2oq0kQxAG
cP6RV7LRQDGWraYaISRqHfaIWc/DrEGyBdxzUC488MkFs2Zxp385MD77DkEv4skT
iroblaUNZc691aOI88ClQXciiVEyo8ZI1ybtM1o6O4aGQsQZoeB3HAHsFRQI5xLa
aYlZNFNVtpaOhATzC3h95GtadoO/1n9pPF/BbpoOn2+gNt3llDMWFZj7KU3iT7KL
6ZPq2MEOG2h/ORb9l/D2CSahD21hczYmbxD2bm79BfN6PLnQ3ivgkSmHwC2cYUSQ
5X8lRrINMJx+W8aK6VgRRYBJrLOhVrciGT8BQ8b8CLgARV3qpTlfmzq7rWgPYGyu
8ovlMC1nhKPJLKJ1vHYkxQxB3+0f0tQ+5QH8Ff2iaZOyx/IKQ7k5v4E9HQF5HiDs
7zdSf9fOV/rkqToRqxm9FOue2kQ8zSJixGztguoXK9bDfr0rFLfvYKVODAJN/EjL
kqjh1sZAxN3Z6vQyY4XGrsP1Ov/4qz4ZA8GT57z1W9ywPItPbacPo9DCH8JtYRFt
uAsAW9AN/aYxqEs1VLbywEQOOQu0OzEvY0txdzuiVXLUAm2O+Cpp3vwvBPdZc37E
nEzUzNQhr9vM2XKB24W1usiiZnPqKzDt5+ovjyFp/NXPpLHzlPBvoennY3SZdDgs
1Y5G08OygVDKUURJsmeXTW2UZBqXqLvnODC3yNduSrDGVa/sOc8iNknYDJu6Vgf8
E2qQbGLnJ+bWDicoPy2syKD8NQDqjNdbetwV51sw8wAYL8LP6uUjR+sOeTCW8Xow
ww/6e7twQj/H8bMrdfDHfas5Zvcv2SNDLKasrdpcqDJ3mLtCBFkQj4rsh9UfPSQu
NjwYEZxnDOojKmRP8nbZepwuva3uP2MF5gL2IChbMuGrSFH8El/Mod9GxJXc4YzJ
2aA5APgYN7O5OHy0n117voj2ULMOe0yvl4yup76n+XVQdkju3XQJ0Ri/xWGM7gD8
NMvQbaDU/gOFlpknNyTY5j0ExlLDkkjZuLwWO/LXoFDmOE9OwDdzfMj7tgbpb0Ek
Co/bYkJRt3QXt0OteJFqosf/BM0fDBDqhiy7VcW6Dih8fkdNX1cSJBDlbrimXeSo
1BQAeBqi4xJZKrdcLMD1N66pPQ8OgLrMmmxurQGA8EXNi8RLrPjMR8n630lAoaTh
NXtbXDMPX3fNdqSRY7AEV3UmMb2FSFreVL8XNy2G3Bf1v+Yl8mjjOFO2U0l6K1SR
V5PFCTpyNeUEgeGlsvoOmyLR7MNXNmqVK8kWR08QOqyoq9VfAfgJF01HyjOhh7eg
ARsatVn7CDvuwpdU4ecDzfnQZShwX3YotyCIbfV/8iA0E8JEIyIiXZ0skgkZJpDp
oMCUQOKEXC/2MTbQOp3WBvnHtx1IksM2m4PpgOyqAgo6lhA+gyeCHT98n0xIXyf+
j1x4d0QvPFNK/MEP/qgFHWYO1yjt+Y4Q2fU8C+qggkj+wWsMW8giJhFR326m9igh
Gp8ecDyq88bTiNvDWaF889BjFuJxMhCzx3EOHaXDrGhQrzPIN/TnMtlSGyTO9/Sc
WwSovV0zxutKuujklfEHJQa8f1rCe5+E07EPV7UTFM9/uAqOK7lxy+g6h2phKCxi
yg9a00xf5o3mMsuvUYV6XATPrtKRMkhT/nu1ldD97eD7zldi/5jrdGJQC45UuoQG
B/r6FAOH47pNIk0mTg9Y1lKDPRo3RiZd/pdmIsOluzcN3eYlsOLZBvhl9/ZXZEXU
EdQuYe21ILt4qPdoWdK9Mfax7lXfE+DV0B5zcCu3sapEElFEpL+ir3J87B8471Ll
ANn3Iwq5TaSAQxqEV5NqRLQLrEzeIutb7rd/N9GX/4mNQ40+wImkhZfQtx1Z9T6A
dOaAT4e3OQMLhjBQHR7EXW1eU3DMJKnYshAVmhvwqfDvzaaAi8j80cIZOwlf4ddP
eK+ePxjyTTxqHRDTS82zqPRjOnt0atus2U1aTKjHiQguTwkfTunA+D0Pt7BWZT7r
74mpX6yzukBHkl4eaMkRLm/qLRA8WkxoTJBZ64G8lNffiUL8pZZKpSl6D6vEc1pa
fwY5+eAdX3ofPPnPtY+1EfXQ4KJ5QjS7ezNyQCTxfWtpR7PLUm3Nvk5+nusxvK2/
biTY080syG+PKjCMrauUOuZLNCJQfTa5zFWMLeoHr7SzFj2tpRJVWraY7UFKOjZk
zn3ZcSgCl9te911NETQfBFFHkn4prMf1I4Rh2PjKMsUFOu1ceFCJEDEQafWEOaMs
az2m1bTvFDxsxhVhtkCE7Eq89w5X+sLnCDH1yz8nuNnsPzWTr+5oExHhVZkbAiKd
k5dTsY+nrTPNDsqhxTgQPIrR47DR4cVzTQ1AVsFVJfLSTijPdxQljkBeYlC1rXIG
9rEI9ACq/2cetTY2vdWnv4jvarTTxV0Pfjy3RQ6/hf2Z5lXNZZkNnyPbSmIUSUl2
knpi4saVf9gpzqjDvTCwio5e/dUkMwr2/AYEo5BKmIzvep0fkINJkH7SKm7izAZP
hiwjhCAUCwIVvGhGF9pmTXYL1KvyidbjIp87SjTubYSRrJaCQsr3Dp1/kDPX26Ef
fWJMUMz7PD2MQHDdksA4IGZ4so8UC9kfwo7u0uINfxvo0W2OVc2X8fobZBhqi+FY
czqCnvjmk/SyQIqjmdInfhK2+paXeltdLgxaM1TONJkksXMH5Y1O87MGoP3yVFLK
+1Iq2jTHnghd+DqHrKjYFgGZvLz8a248MpsVAcOBx2ikpaEbzCy4C7ShTvkiZ//J
0I1xTK7rl9vVGYcvOrOPZX1bwcmzGTMVB5f1nC3sm5uNigAbJGdPgq0FWHPuT/vs
GsljlQKO889WIZbBTsEcd0RdXvrWphDElIPKdixFmT5LLPaC6Rtcd/qWeRtb17M2
jdu1y36obvutWEmn+pezByZLcqwijkAdmtU4LJbIg0aLMtKlC8DGKz9FTS3+sNEg
Gp4O4QbPwYUQGRkST7fRff0WL51mP0TkCeQ7zdHBdJgAPnRyo68IDjzBqVLIZXyb
a21cEUUoO/GJpCDsOTF7FwQJYyWkFbHaTAZe3ALVqDjuNR3uTei5hAKiNveR1nEg
wuMlzkoEHytDLysU7Nt6S1uDUnHJGT4g/w/hniP3YqCWnA2P/ldHFd5MHOB7vJSs
LKhCHy2KoLtzST5LnnbXxoQ7g/XX8LOroIWI+nBow2wq2caBZONwLRyuG6Mgkkef
yiRdVIugEchY4cBezX0pajVo5mTeiyR/MOwbmGfDycM1P5SQ7AH0DFnmW4r0a/IR
TSEkgrWD7DCxWPZ718XzKPVVP+jsD5rh8NoMh88JlLbAQ3BEzt5Upso5Q606iPky
5ujp5c7m3LCrGBO9f0ekvi4ocq5aM995gmzr0sgcD8FKFH9fLaimhlepUGqw9684
bymwUhJ41fs21FnSnAj1ynzo20dues2+jnDqbHC7O8jH9ab3+vv6FABawGhX3FVf
EPzcdniGA6Yhpn8KD6ooRtdFuXVkPd0IRGArrhLkDIzWNjtYtbnCumM7G95LCHyT
aPjKmNCWoHqq3E+vX8UlC7ZProyR9EFUjvz58Xt/pVfihnXoIQglcR2rSyu0swjy
OcaaPpmIxoMV0Pjxck6iiqKqWX9TUPYeNhnqQGzjy6gDCMCY4GROZeCbzIzmW1J8
ZNiYFkMMj+Ni4CyPbTPGSb1TmpX1IW96tw3J3JmwbXoY+bmNoKjIyXt4UEFBtVmz
8c/ks4eUjgaNlFFn8zIpr7Wg6I7n/Ik2oiXSHEExQ/wxErIhNCDIwFJcLP65sGQk
9JMfJ6isIGgv5/p5cPsCNJCZSTn7UaKwVmpjPGXtQXxAZnUmsFR1/3K9qJZ0n355
6ePJ0hEwpqn5K9tBjdMJSzWTwC8WqqIFFKhQib08xge8pMO9AeAIfODI+DmcS/vQ
GBExXn7hvh6BrHJdppDsHWP55z8aItoIK4UZ+8CJ/SuxdpdHSP5f2j8E8AgezMqj
0Kvt2JKpqtcg/iBJGueVoyBbDQjGDqLvRTULKmfBUdfq/kOq1OGfbjuuBvGFKBf7
41fI2oPk20JPK/EMWW9FLJ1OdkFpc8tjRf8mW2VMCNtmfVi/srBzBNuRm4QX1dyD
or5u6ODYrThtWk8IIKld77LdYPieNf2CgfI1Yygv/Hoyg7dq5pq+xqA197p64xLB
niaskfc1JiZPLD1VuigVqNmrIy6Ialm5FQcPUcFJsD6zZc8Wnh3lSIjsdlw7GK+r
gCbtDY624RMuq9g2SBG7990D3+xwpPRLSJs+PdZZ0eDf2W4/d///npwxs9AVsbNJ
hkK5IX76CY1HkWwSpe3PworP0nFsGt6MFfcW8+SxJ5UucHVj5zjup/F+733PlSow
DRPTL+JXemEkITkIjYya+r1G5qF4Buju8o+zwpp0jOUh8AOAQhPgK3j6zHEIddYz
9JMN0ASLatzHkeo1R9mgFcMUcLVncQrSRFNsfzA+c1JKoOB7Nivk9ax11ota50oR
W0Can+M1hZYCryp1aWrfl0ZiwGbFDqVODxQbKed2k9hgRddVEMFlCASp2NKUbeAL
uEQwys5cVgO4zKaDuHcq4ceazVrY+W2hRwN3xmiTZLMlzatTeYV6jXLLeWLryEuB
e9b2oydy6TlLDj0tlizF4vpHXoT8hUTD02dzVRnRPOAcJNmzpLVB+GVERa6Vbyc2
sQ0xWAQS+FNXdGaT3cqFtIzM+en1xAiPVX+BQZdvjeXid6yhjk2vUMD1z1qTJpc7
FkKNfruFqPCasGpfMgdl8GqTfnz0nTky7aUYVw6XZmjIc9PZZJVBdI20NDbE/lhY
nT9u2QV/r7/aFuO3LNzcodcRItZ8yVBaFYjeB5CV7Z3oBRV9hxvKBvHdcI8IuClS
9zIQm6BZTJOJDlCWDccm8Q5mDdxrURG80Gr4yvIhc5rLKOLp+oZvA3OXD0SrC5C5
cuR1LZ61im9YxkiUvhwVJ0z8JCtb6Im9MKUR7LC8qunNe5kChNwD/BqM0lSwGghS
V3eYVMIiE0i1Y+UqubRaQAyyBA5XKo0BMeYXw/jemIEo3PoNu9nwADWphZwf8aN5
wREznwElkQyDkMWQfsGnyASf0sauLolBJVhpFOLk2JAO39uzX2Sc2zIQpH1bWFEX
wYKV6MrdoEOB2VAPNXfZuFuWtjY2uBGpMqTrreL/fTGmtrAQdMh7mNRQUMyWWFH0
7m1kr20ixd4RszkeyO58hjqx6E7ZiMXWJw/Eyto+eXd69blrITvn9lfk/CCaHajr
9p/WykSblFUUpeNB0ZYp8ikrp2GJdGtT/zgoZB7UOZs0dHFHOdysYvH4PrG2tsEw
jPry+cXcwJFGcrOhD6mkVb+xAxXYkuBbIjXv1/q52c55WzIQ4CGaXIRcAsYzla8+
oDN34JNaUdjFwFUEOx85dITMZ4r2SBliHu6LVENO+Xj+n5SwGT9DFaG9/8tkdkw9
JS1j+HPilIooD57NYcH2sIO6ycjizdH7jRvXJfHWSOvyIOORzFO/PeK+m2G2Un79
ApFuhHJYsLwV4rNvfDyeCq2tHNtMg5NmT7RBbuiDVIkkVihkDnNv4ekcW7blMeEb
JFwzBco+l0uU7q24OpHu8qSpIDg3RNP09wBzCIPd6UzHiANABPY8rDWdC6QtwVOD
k7/ImbMzgwJGX+GiRPGh5k09Z/jjR5jiVslK9FIa9F/uYQqtiMgUQ8eeYO2M28/q
Fjbt/MKzcCHyQUULGTKRFn/TbAUZD6Airs0iGb5GoZx2u3UNhwKadu/zosmP71pa
EcdWbsRk6Ft8T7ozlmPOG2BWjHSgwgiYmUr6jS3lQL/ap2SqaT70uBbH2Y2J3aa2
8Vu7QIJGRxCEl7pLINpX0TiwOgAg+9uhJWJB+euPDxGY4rlPb1HpH6DzXv8nyexH
iupgukic2FModJQ2fLd5AheAZ6YsnvXI26rzjmbZjdcwrtsx8/H3Qs/llb++NBzl
wgD/3wFlZs3ASf809HG6Bur0w9dYh/Z+D32FWeRs3EAYkJkw5i34Ha7n0tQH3F0Z
JxZpe4enrbr2+jV2xoB/6N2JllH5QMRiq32HsweFfUZy0KCvurPm9b+H4rwNhh7z
tURgBF8BIn5IOyIV1G9QMktC7tdvKH29FWYKTg0rA16TdKuGV4FOJRorxD6hlxzJ
h1xJTDYrdtNufKDcRhbKFXZhhl0BA0vWkblNtpaDHd4v1PCnY8PucAfMVray/sLQ
j/PXZnH309nRiqf8OfsXkDQbDsSxUCXLP4FW67I4kmFY5vTxG9tJk5oj7sN1AkSO
gDBigOuZLokHX826Vxx66g2LoDlqHZdeiFqCFVFlfvWtHarpcpUr7NtP6Uc8g1p2
qu1vNrlpVaJhRNaH8nrPeamKzsehhRojO5Fg/oF8ea4S8RWIYNTnvqKY5Yrt6ZOz
Q8iuNk9JkosRvQ8e/D9z6dTlLKWBJOvzzmErZEwikpENTsJPPsFfU38jI/5k9YGY
uIBCZsOKvP3lPiE6f/8/pJLumpLrWR1yYyuaShIvJq5EPOHXA2ZvAZdRtfYn8P48
cWJKPIubIueHOe5MJ/9Z9e4Mh3OLcGrLSkCMR3smR46k15WPjcI7nIgnQ7h6OW0L
vfpWc0np+r2j+22gCCbTuocg/w4hGSLcAjnWBlV1Q/XZyxrNddUr64XoND4IToy1
ukiskt3FxEg9AUOx0pkahf/gzhxC5sMCEcTANfazYqXi/vo/5UEKj+2fJTEq9zmT
QXwxY7S3O++hdB/82eBZACFCstPvWYqPLsjOZCgl7Tmj8o2MC3+mn+1FFR0nWaID
Mmx83dy+lrSdS2cg7m3vYFC/DYCEjtXex4SqznQno3/hNbMXY66P09fbbAgMMRWY
dus0u/kPuHVTbC9X8HdU8C6GV+ri7yQVJqWx3uLO5I9T16YgXGXvqQ5qfSbHLa1z
KHF3HCcTZorwhoN99Y4gHqjtwcdx/jAff2kzSnAXOLe/EAWNffZwxHIjZbZTaGHO
+Fhh3Omd70d7/ig/bfC9O/fqSn8eeNGyEZHQsmrlGcA933gr2cskFxD+Yi+/sJHw
SsajVNmzPBfP0Dn/C5jZAy1uXStqvJTEplQblYidJbgG76b4xax7hwKTvGxpqQ/C
spGAd6PeE2dBHLiZYuqXxhhWG0zQeCuvx77eyT3CLCtNb2viIJHt0p7x9ISrITr2
9R2dMLOekNm6c9vJkTPLpuJfjn6r91sapqr++7TqnHrBznxnvoa+POqVbH1zdqOd
uF6wL+aJorprusBlZqVQv3rJAgi9dN/gZX7CGfZsIUKjXzMyhl/aBmlMf7SEiwdt
GpvmNRZCbyf2PrMxb4uUTDodwPhUjAdpeQtBPNfRYqfa8hO1U+azYeYGlPr18oZz
1SliHi3KDzyLimQA3qhx2Dm1HB+wzb3BRpE2QANHqu1IOjvmv2sHsCsMhT2UnMRR
TW85MgY2Rdnbyg4Jc3Odi9QnDvNYux+FSsd+t2hz0QT7wf6iC0/SC6qxJAJ8s9nM
F+YARQdeK7Bc7NP5pag/vRU7fi9U635bDHFWayz8MxAIYvajzLuVx2kAlR5f7Fdh
/8WAvTmy6U/18YJN35CCTafWCy2X4N+DWJw5KaA/qoWADStu7RwBRxQdLjW04uKr
C3csDCsrkQOU3R/iolIcKAgT8/ujzdGVgGMNt9Lml/J26X4NWLerCAuxO2FCjus8
2mt0H/BwgsUF9qiYgoUo5H5ZnB4c1lNd86uEzZAplFW+3owcYOx9HnmYB/R8CpU8
+xJSIseTkOM1KgkH9z/aVF2ZOqvjRr+nMWkZ6FDh++3somIkEfgH9jsOinmzGdaJ
540fR8xO7k80BWDEyRECh5zO3v3FxfpawTmFDmUad56lJ8VsdPd9ia6Y7hLYQsU0
IbU8K2qxAb/NRTDfqbQxZOxcCasudUkc4MHaNN2FLXNZdKrupGXYQF96g0pK+NcN
pna47UJEcDU3tyek59LlKuU26heLHJeKHc8bYdy/HOSv+1+b9tvX6sbeMN0Ek/LD
Y0AGhZoOtjIX/7Bs8YIwEq5WdM8xkkTcOhzFssLLeDne1lXlL0OdpMeqm8NJAhc0
3zTfTz3jjOJk6FZmGJ/PjBGEPUDpwJMsmugCVHJtvtn/+QSDnDN0Pq71AoJReCRf
EKuwXVQi74G8wHTRwBDhQNAvRdXoqsvDNjgfp73WqM1T2qRCYCEi5IQ/BUTzClls
wFaERv61XJ9Z7oEP3P48VkeVu+tm8NNOPGWFi6R0KWYeSbId2njuzg+GgUrCrR9S
6PUt3bLD/OtmVx4ybwvMkV7Fq16rmg1KEEtMt1ogxn7S4l4iNUBHVDVDoa3I1OZa
NAJ4v4MPt3tBqgmEK6ObfNke7dD319WVsg8tetHN1hMW2KD7aTIDqX2yqahF7sFq
ovexrLktgyg7nZSvNay6//yhS5eua7OUEFrwU3EkAXOlL45+riRi3Hnej1gZNyww
Yvbwcy7S2CNyOgr7tJ/KDaySrY6YFUH/irhnSSxto4o3oX6ILcBxNl+mM4vcdHiO
+3+0A0sf5qLXWqcc6EUnz9zC1Fsvn3d+nWmgIAmKDMnEoYjx4v+v0nDfzcLejfx9
q901SNxuw/j8MKAwOFp2g6jc7Df40RPzrWfC+Abyohn5ZuS+06J9i+iFmNo69A2M
5mgKPg8KkTxR5WpAZQ7sSH0yQC4+4gVQjggwvF0m95/FM5VoK4aZvH3Z5Hs4XWuN
ZWL4+c14jGjfT1+Av1WiKCQRgzP8jnh+MvkN2AcBp9Xk6NMy731B/M+Kdcc7mzta
ZHq4N6onecwrk/IXZXgDHtrJrsIZxxZ2kMVHW2r4ZAZqqS22pZNIRLKu2I7GGybX
7L8RHXg/5N6Qu2NEaiudOBDZIfsBDK47a/SxA+zyhIBb9bt0RNUqejmLvwWQKE9H
awxeGOCpqzzKqFQWEaoTL7iuLLUfe+feW3RtlS17GgdMbsfxiKyT0qb/0FNtjF90
vR+m1EHGrf3w1lFPvCZweus5iGt9ZkmBUCgsMPughSsVQj1GJJorNNl/rvB3OX8m
9BNpaSysuWinqof0jZFvQ4UvCqMRpvuKxKhzpbKVdpOyNwYJgW/2sFPko9yrno+k
676uLyQYoeggz7/9BLCdxu7sQW8hmf2hJX2xCEzkrAldwT8mQnCgUd5agmkJcNsz
BekKCNGCrZbDgVlbq38+KZU7DP45dy50FP6Wlvj0egXT7hTzG7lgxqJ05kZuUpcm
ZHWBJutAnffu84G6xWQSkRI/ufwbvphWkNaiuMzR8QroE98GeFqLL5SLnyHt0mRZ
/FqO4SJwMYDtYMIOBCtoIaRwyXV09ZAmCfdzDnOgtAYjIID999053s7cwbNvDnCZ
uTy8dF1EQlTaPvZqkSrC4ynuAt8XX7L1ezAKYH7waBMa7y+Jb92Ng5Z6YbSTGZ2x
L4iSPDSmaDuNdNuHsZHStQVrQqdAQ+AQREcyb76pv5RZGVraOWZaxUnEh57X5wh4
j6zcpm1hpiUOPMxpabZ5Q7/8XXxOTDOV6K4Nte/tqiwK7KuokYnkGy06uKhB3dYe
RPhkS9X9Jz6Ybnp+n7hsE7hoVhFeDhVy0CdUkHKGnrQ5tuddu9qfQLaqooJICrZ1
J3S9IPoyaKNfcM0gnfNZfnFmFx4fwsMziLu0auH7ENmGccm18qk5RMxgLVEm1qDf
XUI1YPfKfv2btwbLV3WxVCEMhhEP7KwIglLnircArKDoYjFEHAQA3hUYput6p7hf
C78vOy5o5s96104eAehXzNROJIqqQ05GNRLO8+1mb36/zr/oykTC3/FYbdk1Wca5
v+EBAsYF1kMNm+kP8o2sLvgSKxg4hbK3qUAU3ZcQLrY1+dGroScN5M5oIUxe1RCq
ZwR07KHjJ8ox/3izydohTPxjhvqhmUi6YrMESbHbH4eFllCc6Q2Aia2RxQ3G8SXA
4bpMhFaD9kFvXhL0LQPp5A6+5t2PIvPaSRfO9lIZJGrXEyWzWECjqbYQFCqJQiKB
8cWLRkM7Az/1gYM/Tw+IsM42daRjLLjnAonzGfYR8a9PDEe2oweJJZuc51cSL7Pm
ri6UIro+8VP3/kmcYPDvrbEYPndsUOAPoncRKa2Do8Xdl68nyjT3b9soJE3e86/O
j0k1GZxU8CveC6hVVnP9Gqoay07qIsxij6EvXKLRva2R7s1ziWG3/ilHku+GGThH
eekpAGhXrm1GQwtH3kp7RhRdYmeTTn02bIPqzVMgnRBGPMzsHEr9WFpkydxg1ugF
3Jk1tl3rs9DFCa6yokvYA5IFGF3pqJfUc1yqBeWh9lVT6NnEfcZZsyRw8gNsqO4b
vJko5GQiqTsgnvvACQZ7v/iJB2iAffRuPPXgcZGRm71Pd5+TujibNqjicNlyfEys
Bzzj9DBrRrgOkKZef5BpfBmGX/coNMo9nDlEUGhiGtyoXHPj2DCwt6Z9wLu5GCqU
/43lWB56bobuEQDsCzSTkZOAeB/biA0HzQeZlKEQtvno3+R0Qf5D4nnRwM65G4u/
Zl7Zyhgevof/J3xhTAXPUBmppaXCP0e5e8utMrNmz7qBENunI6nlBgrYUnmd5yXo
4igstKBpvif4vFYbbY94pAThQg+sR9O3yhRbrFY2Nj2AIaeTfM7q4RUGVgUK99q0
wM0fcxuZEg3wuXqqBwWrvLOtsS5XiLUBw7KWUOIxgq1yiR/E7k1Y/ON/27tvmxFB
49K1zb1herHkF1gNyf1elJ45duzAzTJ1FLbIAdBw5dOhTeYz517jMSrhg83xIhkW
FQ+rGEVey7zXYr5XDPPCv+NdNMxgJvt1AT4zu/IwAk8y8dNlbVJQoKrjonMnOrOv
icnB52H5y6qd7vDfxh/ntU8W8EfU7+74Sti2IE1aAwWrnrfSGMwn3Noj8TuMT25/
Wp9UXRxUo3CZr8Ol3iLskdqMNSlv6KIURFlmbV0vMVOo8L5oWht72XpJr2cHeWHl
KHt98mpuLnMpJ+TwgE1FJhXmy9Gkz97BQwpr+2iLf3+uAv4o6I8TV3Vaw29N3yJE
j0BCAuDipiwFa5XgnYx5ZHxQpKuy0shW3hl7ws+QjqDhb65BBHGUePMpB5K8mNbt
3wEjVYsQXuzGCWaR7jYHqdWiP0JI3eraEacTLSuOCMLOq0PAiqF+rcoRYPJhVYiT
DXbVCRFfcEMCtkh/mfVVsjR/GLIC7+egBvVYlLOWeU+KzJ9diLaGGYb5cJscA6/b
6mIjSqRjpfQu+gsydSrHgokAFQJF8PyhRNk6+hGNZB6sJB89cHiwxCpHWQhEFzAA
BenUW5ZWX0FgOGzYgBGctutNQQoqpt3E7miH9G9rynBwkZIlrzmt0yS/P4W4lF67
6UCTHw4GYm8RPRvAB2/YweGMHmclY+zswbhEjnrSIELhEnpfVGrOOn/9Drj651Hd
ea3H0mioScg6IDWBCQjZ8+12My0gNWNwMMYEufKByIGPgiDgO27q48bNEfj+C7RT
W2fRCFClvh0E2WHeFX/UBuf56pRe97dtEYaBxmjyQjjd+t7isYwFKUtOhWSmZUQL
+TRr+oovsoOJP6d9E8eLA49ZKdm9dcm0sfT6PdlFHpAM1rdZKYeprEjFRqCD5S64
IfA/hjCjqXQxYQiHo2cNbnUNw4VatSDJdJP4+vlSNllwE6a66YyEqbtWAs0sFC2v
4AV463NQIBbtLmam0VRC0qN81AbxjM/vd7riOTjCBS/4hODxNNTvIJ3lkpcYoNlM
sIIiYkop9e0zmsKJe3B0aUdkKi9hxlhg74AytWgycoHAeifcK1Y+2CPUFgePmQmw
s1QJVi0smcLNukvu1qMsaTL7kF4bXHq9iDZ2XvxFEj/psZKGPxvt0rU25l/CXYQc
Vv0wgP7q3WjePUzA+U7Kzg5Yq9v5SwQoWvb+TqRVt2EBxmrbHP+uoDVIauw7byEO
T5cJVFqliQttHimaE/t3c33ZGRtC56HlojCmyv0v8wjc7EPbwnN9swlk/zD2qLhY
r2hHdDP27Vkx7lFJe7hxyzYPBtTcMt1sbsdUzmyICxMpntHLzT18h0sGdXBxdi/d
IjSrxQ/SDi0fgm6DlMcqTXa4M8C7nIVN3/iXckc9b9lSf+9CYR3/I3XuXcA8pRO7
cn/QlFRZoSnqY7g+v7KDN6l/40bwIYnjgY568zpbp1k+ZAEjm+BhzvzTM8XcpnvE
9XbESb329cjghwKEIZtk+sTWAlpuCQEQVCzX5Lh2QYXV05umh4tY50dhrdbGoBli
rZ8W8NejuMnPFJY3bANfwO3goKFwsPflg0daaqANkTt4GZwXmXqfS8gpxJqNEQDi
JDsO/mYirrErZ2/PwUuAY8UTLNCsbWadnA02q9cId8djsehyfgSxkMeXxAPlJAyn
t0mZHw7uZStFeaEJ9ipXx/6+Cah4BVn/6AXKhMTeioAd6MtDEXYban9vCTtIGjad
Qei60lRnp4kVMM/UjACJeUz8E2TBsI/2o7a8ECGlJrR8zEgotm3uKe9kybuxCpxI
U0A02eFJQ8QRp1aGnSqgZi1RtsJOTfSoN6iHb6zinzvJgCDLPPOVm2kQnB5XOxJZ
76B1Wqwo7vOz88X08Y/Ig7ydNwdWCAVZGoBc0uV4Lh91LZ0ueQQyA7+O09gybGMs
tPT9I90UoxpqaBwXUSF9aiwKvOsFchVG5q4j+90JbsWNWF4rK5K+e6qHFe2jzRyv
1y4XJOCR+2VBuNJVPds8XHkVkQp/YdrYabh1SyQcbPjxII5L6WyUTutiJaeE0Tf1
oiLGY4BQzeRR98am0t5Fwoc/t3PGBPeDWQryISeyURocF+Ue3cf/c0rJK3t17mIp
Bp+lDz8E8BqPViJxu8sk6J8fBpL4TY2QK9d3t1AtQiSXk/tGLroq0X4Kt3mgBmLT
/v3Yd22gTpI38Luvgp8gbMAjDFzgEZeO8LDluVfvLUQKoeZuBi79vBYCPnt2ZIET
XhBQpvfjGWW7m9KSq4aMG/YaP23DYGY99PqEmucvSK/et8g3mytpDoVUL264wQ/4
QdHB6uDIezdKG/Aufq+mNUaoCCAqUVzpJJBa1VcEUp1FHgjpN3FPJGKOaMwMoVdL
1eIpqZAtJOhBqgjCXobnsgtn7FbU4bMajJLSuKfkfr/Nh8jSHAzMcFdjQ/NjG2pW
Ach6CIwKsM0Dvjjn31p01Y06qFH7kMhLpWyb/kwZzpqI4goThf/pMn/IFC6LAgX2
shAQOPJAmQc9ZMnyMAuBaU193udJrXSLEc/kO6N9YBJ9DX4vC/R5Bc4P0q/yxPHw
82tFaz9OK25OWydNHChLxR1CCoNV3rDgzlkxrUBLs4jPJ5j4q55l3WUzUXSn7JNj
g6anxkwb2uopfgKsDXj6xz3InkB+ij3aMei8xlgxeQgolkYO/jSVbhvlUm5A4eer
OBwY09K21JFoXrFjEgz+Ker4IrXseeya1d8ZRZ7PFmvgI3HAGU2NUMitJ8t2WzKb
C5RFZ6/XNjc25OXeSRpOXYye0fHGjvUGyrcZqn7AufAhwOK7bEDQkdgWZQihAgg/
yH69HbUyUfGUKy6oW8c26hv7pZQ0q1nn+SbNHK0gav6rSSgL8e5z0F/6VA7CEBTt
rM8qczMwLL+Kz+cWDFwCwSoFxeGY/cyB7swxjH1RsMBuv+IBfyUfvOY+W6d9nMxF
qr5/jU7KagvY03Tj7zWnz9HbDh2IzPbiJFRviQwjvP30BiTPMoYuIggQOyQZrf2g
mfBnj0ac4dMRd1IYaqpThu6YLa3hGlhytHvheM00+cXG3LDcd83rmzQELUj7g5ZW
ypbNmmytYpin+V3II7+nnpvyiwFiEeSH8uMXB68UOVTEDJ5ZqmfS8dW7qwJ7o+q6
4TWKPcjCA3ozu8KKF7RBonwNL+kUECWnA8IyhtBgyJDG9v1JJ+T7iCbxcFndYpLY
cysmmnsU7DOGOwbL/EPjMQNIv07VVUNYVIdoxKDXuyU2E7qXcOYzLA0NaCmAwW6J
WCpRRqs22i3X0XYbeNFtlx6VNdchXk2390mnuDSQb6gFK23dEJSKxHEQ+/WFgMdX
wy11B+rONjvmScpVeDoMY2fU7z9iseiSKSPzpGhnS6LScTAnLUUSpnxRcblr/3Ov
N+cCOjCnKkU0RAAyBBaMyPiaKp0ovnwpjsxTZZNDS3gULL5BVr0+WXtSpARWfrYY
9ObUPKcHdwXDQHDEHVdNuYbIJUJw6XmaWrUY7YBS5AGU99QzI+z/lwt0SccARZe4
i+IxiHARv7lH7JzL+CagdY5vfLAYcasKSwPz07B0T1z520RtEFKV455sgtOlYmrc
eU0YzjSPAdWP3Gg47dg0dVhf7HhHWO+NsdxeSwekwc0PVbwJswzEV0Cjbq3ZUIRT
1aiHREXSlyBr6KDvskPC9Vb1QcenoDqLkk9ylaA6RBnU25iCMh0mswdcAY4Ev5TO
GXxkttogA6vLw18g2KEDLOgI3RuKBywLeaO8UxVq5iLsjoxeWrFZwU8L7FhJWCz1
rZXntnzewNhVP1DEC0mlf/1uT+U718d0O0wsKH3+5/2p6iStnOkeCgkw1EuVHH8+
oMGNtxMpfg5h1k4FqWmdwQdEKBQamvGl/7v4aKAULl9nZr8XDQd0L28C6qGSAVdA
9DWiwwAwgkhIhIMxKbeyld3F2Rpe3NRXyels2lt9nWyIcKHJDr1NxYdW+uVLw5c4
ZLADl/8g1dabP8NoTh+IZobTL6Vb2YHPpEGNxFLr6wyaGpRYYE4i7x3c7jZ5BUA/
AtOGQw1rEKNPcx+vUnFey9zCuSi458XVSZegayJZ3mkjAbsWm6WwJ1JllVjbYGcT
Ai/1nM/EamUdtXLODi2Zo3nu1VJznoTmRmvblyXeJogr266XnHzpnT9/VyAPb/re
tKLJOG3XtUvUgbzLr9eqp1FtOMNeeTA9R/uxqggVOjcCxkyzIHOM3O0MI+vQEjah
HrqqLXU6Xw0vjEZo9bfGf57z32Be8uHJe9SRKG7pxW+AtgzjRekVq37DQ1IxY4JI
AlCyXUHdZPZc195rMa20dbMaqGVF6IRuDWUDGZuDt80AOmdMxBRk0lLQ9svZKP4j
rAlRDkjxq5xcdqAYwZXvvIeOxBNSLUxgyXtnshYxbvoZNBRS5j9MpOtQUyE1A9Ey
wd5yhYIHuZVNtS3ZZALZRwtRjCzCO3k0K7crn31eXqy+QWoBMS1uCLn0hf63EGkE
HTmOL4kyGf8NUEopHbZRSThwwOGB9aU1VcXA4nmX9MaF0/BnOr2HV1jE8qLGU8Re
fAHReWiRyB39XkmP2+byLen/tl3MMgTFb+FMAuV+FG/82Z39VwF/yZ5Q6Mb/B45v
K3VCxqlEFhLy0r043pIbah5EHNDEoryORbEG2F9xyQvELVajkMB0px2xzRd/3q3S
2c281uWpECbFlWKM4v4wInFzh2rqV+69F4MLWW6FW7XF/5wwCMpPDYUEIvJTd2GL
Pb3h9DDEpWF28FfbI2jndyvOeRnf03+inm+/JlZascjdbYAfFZziRPk3VV9+x7E7
a6ORWzNPqOxaW1G64+4FgH0FOc6sm5z0eJ96yvHSpg7AmldOZTlr+b7AUqqC/nlp
9A456i8puFPNiLSefaicQvpRzpdHgcon4SRf2k46+3NgvGALP9sxmdtqo2TW1+Hy
whH/esjmUzbI26zNpfK2x/7PgTD0xsHgYkPdfx/VG4D4mBPndahut/oYY8CeDVd/
VUfpzkwKfSC8iaMAvx2jBabGxEh1fvtSEJAaMBTnkeHAdmyjGwplAotfuWC/VMrG
Usf6d5VYZl14SoA8G7IbL462yXee8UVOuwvJ4pbIRK/1q8RfWLzdFm6rvyP321ET
4AWPi3oGRJD2BeQRNKU1/MrWopKmBeB1Ohkdd9RkZ0IioSL7651NdiVABIXU2nQ4
HZ8SBGhXJtPkbeVWW9+g0XNTvPg+u9S7SIuYsQyDpgMLjMfhHqmosyrPd/5zeGMF
hf30IZD5ZqSqUdBekVABcJirUvw1+GfMplNkPbLTttnJoWATGZWqSQPzcNZe7uOf
2SU0IQpCSSDbi6Au3+xk6f1sAwZB7nBC+f467B7oWYjsC/lCkzVs4M0qP2nl49X7
VRhENQzmGOsNGMzheSHJRTZPASlQl+D8U2Gt0gWqs4N8KyFXrBGDS717o8DbpBpl
gzQLF8/g8y0ly20iomeZRnrOiWIngSsrMmqsFuf/EPMgTzEyFCPAMJAY1c2peflf
7jNuvqIrGmch+FzXfpikRSefAr/P6pC/AWsGlPV0MWfxt0OFWXcNTVAHOurCThea
cCVmBcntC2ALK+Z+XrVCuHnIa2FJwEWJkKd4lkmkvAPaJ7yWgC1bLu0S7bFsluy3
tHv5KuCQyFKlcUh2RFJ3Lii7rsAPyIRzmLhTXmK9DL2SAqfRzebTXmT4Yhf1xe1S
XlKCGVWWftOqhH/txMiaM3yl9Slk5zfXmlWjfr7LeOTOk/TiwMbfbNmT9DSsspDU
p+S9XHSHs13Zh0THxBM+IZ5XKNfAnSNLj/diZgkjBFTzxnr0qNBqGxLQpbqObQBb
2ot15UsuP975pc0LMwrTwjtT07LeQKl3EiC1T66hBdrg3aRoHpJUPjJcLEHWad5V
UWxbVOAdbyhbkhiT/SQ+KcBwyCsnXG+pdc+UWGMB4QFgLc0nJFowtRjxdMoGbHFr
tIv03AIfnrqp7oZS/u7LRIQgN2wZ523yDDSl1/grV9HlGfejOLyVCnc1GZRw2ujT
L+4JuobeNAlJBZhtznJnbAaF+C4kPsF2JHiN6xcj76j/ogSzid3NjAz4nL26pK07
ahBLc5OOKicavWPoeMk/fJ1XJEOu9k79BTuS+fFit2Z1PQ7xY0A3TD1dZGWMtGFF
WbUCIGMmTYSWz9YdvkpR4y/rfzX0oJWEp6AQPxk39ZTebi9ry39ISynY5W6rmdCd
ZJ9IQ7y8+WgM/aN4JiwN1Qb8mDleRtNyCA+Sn1juB2T5zvHN6/QJs0W/5VsSK7MQ
QPqrabEf0KxMHxEOjEdQin5d4lQqutYwMZsNyTncAv81boDp1no6TqiSoOMn+FUJ
+cos5nO7lNzDrGk6ypGoruW6XJqQz3tLNrF7pYzG2r9oyvjKCMWmHqfmQGYC7aqF
18LdNdflOsPjmck4RkYIQh2uPxZ4eFWIHlD4J53w0kmOgwdfqZ2NKVwQ7Ju/bito
2UxI00WXk8lxUnrXI/shjHCeUTR/zLsSVgpvV1sCZPJl8Y2odxu5ftp/g3Dut7Z4
qcav13WZdvG/wr9nRHkhMod+glDuMzS9jPrMqw7JAW7FmejXyWZf/QSDYjCAxRwZ
EMs+Sa1tVHeSUZTfM0Sq2SWLFQnAOFpSp9Zqv3eRwk8lXqg+eDUD7Q7fW6JjQ50m
YB6dCKGpwZAsBHJh8CeH7ZxA/PRrJ5n24XwfygLqoXl1a3Sjkrbpbf7uAFAYhcFQ
ydizTToikCJiXgCdHiEgpgMWmeBAxJV3D40glS6/8YrrOutrybBxr8s7sAV6AQmp
sqxIDKLFVzMClsXw1JF5MW6MhrK1kWdoETkb6JhPCtS7pno+ym0HZB/VR1DnSJEh
a3Zv5SFBjIz31hcaOje45DvO250QozGfR7mmEE3UNwtik8sQ5fgaYkYbAFw+X+VE
ZbbMv7aBtP/3Tmwdfd5SirZCBGPmkneaz8KsCJPsthWkWHcqw4UfzQOUHaBxOhQt
wQUuwbcGhVhHGiDxLPO0CXM7B2p9GSJf2j4x2XOG/iGyT/ZQ8CyAG6vjNtIz8Q8+
cKeFmOI2IOntMJQXp03q+9hJIN+xcD8TkOS1iiKAPvVDODep0nF2GfE/vbIfKN5t
SjO452KdVFfG+lGoBKOql/jtjVskjcsdqSp59kyfms39W6H+++UvTLqsFH5S/dtT
ngm//7lwI5LmUp0czfv9HFoWVt58Gb6/ijEqywmHG0W9Y6YJvrpVT0Sh4NylGLg1
7xbjYOTBDJJgNhYjFiqKsarzzmDqwLBIyt000HZDB7o81HMkGjyoHybXz99ZFMwG
QyYeyeMdvHtvE6GIB0BJIDAeAjT40Wn515Ytsn8o6o7SkrBzyGh8xYkEpz1QPBR+
NYvHuDxEr+bhzH8f2u0D821mJrcfekyjWR50dBRIIcI3uWvA1EbtZW2mT65LQ4HT
b9yEOmMI1kpEwbGOZT6/hU02h93uKOXftPAlvaOWufVhQebxki0OpvhTiYG7mDb6
StWlOIt4/oi1JMmLL575ypatkwKGyE5wEcs78k+RYoXJ15TAa9jkH5fwAsn9AHFf
6GQFbVjuRlIs0oeucciiSUBRyLujbvhEWfxBU4H1Z1O5B5UhisQ4N9GIYoOcRlk0
2E63bhzKmwUJUnNhV2YLUSQ06M25CM13A18WN75Y2W2cc6TVQOnpwatFoDSsUhiD
UJaNOauOtGJpV+j+7hqlnPLZO+AUzfuLOC6g0XMymKV2IT4C6o7BXQmGTR6fPgMZ
uAkklqNm89ql87GIYv1/Hf6r2FBdfouO+daY9YbMx+tZgJadSCNF0EbAFB8nOFeJ
JgN54WzwIp9geIaw+De9Ml2NODpDyPdlwxG7n4wS7twIQ6fZuBsrCUTf2HGmw5wl
vrDMCzkKb5gTag2+Th5bCtUJI2kbPYXGJ7MMRkGNHlIyd/xGFVdo8zW2opS98JYN
Xs9ZTkXHrd4uMeJSwDH8rGU81Iwah8OmAktoSkRw6K/Vq+RD8jlVCP82tHGBF/oT
BGrwkFtqBy2KB9hmJme3Hi/+IxcOXFFIaRRynVUPyV4Hr2XWKs4rDYh3nq2Erzc3
KfV/ecg0/S30s7XuW8d2qKccxjBDK8yedtvotTSoBPphXVXI2G25T/qRaPgj55no
xUCNYpdeGCB7rYXN3z+/0sQPF3VuMAwA2sNL2rmjtj9kner2Vf1AUW2t/Py31ddR
H2OZl+kU+FmLJ0MaShr5NR/GNVBDH1REZoPXXTin83NYgbSawRD3MkR9j/fT4XZt
g0OYptpEcBsuCozJMfM0PWezKEqvEfIHirw3zx/rebYXxMlDWPEnNs+E3hfhv377
3RxudCZ99Ou7ZP3AYgj/84qxoKW7Gxv/tGb61veLLvMgQWIyIYIx6nBOr8OFb9Ji
bVS9vRozMn2GJg8dZg+gLUU2YmkHINIvUjECyKt/f1A+MoNiQ8hWjHQdL5LN1fPb
I0gnWqG+77s9ByDY6vV9K+PchVdHudEjWCVzKnWmjcWrw9FP0QFLiPIGg+PZMjRF
BGTQ1sSgBlv7lpJY9YuaJbjgGOO7KQ3SDBPN/Zt7qCO6cVIKlsyJK1h8v/J80id1
DzmROxN8XY5cYpP815t+/ZRCjifluERSdv3ZqAarZFQVdQV01IQTCW4Em0KYQuSW
TY0mZ3da3WZi6gVpMTrUOSpey/BG/qD1shHt1ev93ilAXME7s9QoqoC3bHdR8Sr7
0o9GaJOdf3Z5FEZFHufwwMVGPrhA7Sif0cRMqzr4ayrVkB5pFmCnw7E9vyKcRF53
u+CQfEgiKA2MuE/PiP+veJM8BCrelxx4EoZa/hH6pCF3vRPbGA4eQ1X1spzFUM+h
8XS0s6PTU1sIS2SDVHZ+bc3zqhzIz/Dy78Nwb7iiMYUACmmiJduFGPEkoF0lhVOX
Isx+iOdWRTAVwmeO48tGdJj+KP5+z7PUbdo23ATY6oiV8gMf+3dQW8gK9bshReJn
qNzaPtdwlSF3eTUbWdOhqvry586Ak/mQPBRiufgG+NHdMepEO50E2iR8k/f3fTj/
YulW+ZFcoiWrwjaHFszF6Gu2tS1HE3EftnKkVxGhwiz8rX5jnwai+mgVz8yBZM84
Vt+33iNA5SswKcflAbbBWdZ1LeuWc3q9xy/T7PSXs9aWulKPxYEACoZmdXUJzaOI
t1/fdQ6JnSTGNN9VdM+NiBXjS9rty3bArr2WJIX/x7X0tDMK4vSYW6vdBkV3poql
iIcltxlYsAzQaEwgMBE6AMqogQD1E52LIYFpososeefRzzlp8NSe4x4mv67m3gB6
0oqOSxo6Dl2eeZDXkrrtnc7n8sTZXPw1eTHGi0N0QXY+bM7iU4Oeo8t3VHoDnifa
h1E6nEDy7AfBqafK2NZbdCZ3l3ae0I8piuqkC1+T6wGe/y8b9K/QGdwy1k2epNW9
u2ESDQPLpMEbXAhx79PSnsnOUrt0Fs8E4UpCfXBnp1nsc79kWv3XiJoNzyNNUdTb
V01VbWFqHih7rUgrMCXMrk1Jqn/0606vT00Ht7u0zSTTr1z8rgftmAqdjF0lTQDV
zzLagaNQOxd3cuj48k+snqcazmUfCrqnuOCpIidlz0V6Nj535fvLYiAWM9K0aJfo
thXOtEaqIdHx7sbT++BAMWekNOQwZCOF2gVt6BMGzFosQs021p0Kh7wxE1tXznnW
RMRVwCfxLxZGMQrAYtz6PHtAxFQMXoqdqZxnyIHnARWB68pwVxq132+iTbwx6AQ5
h7vOtCrkBsKdqVa9XKI7XH3eqTX31pDl9MJxiMn1ldC0XqyLdsjOYVUcPlx00zb5
us8N9SKsvRVJ5E3KkjNllDjtup6CiT8dTm4JTgHi1vS38UYUp65fNqLTrj0RCzhC
dlo6g2N0D4TzFThe2Q5eXvWG9K2Wb/eTpH37RTZSOwDy92wVMm5/ULjMyTzozipU
wzMNk9HCWaiqscPmt9VupyfneYJPZfXpqtURnbSc7zONrgtSArJSjjoqwZmCiUUv
F+qd4ev1lDxgkvtZRDBjLI7xF20tgTtxf1blPbfdnUpdkPSgOIi1JwGenbv3yuFd
nulY6yUaainR0tiCBEoA+06AYpi4FL8FJUq2IzxuLrg4NltricLXS7m7Fqvgmri2
S/x458phZOmtkCuil++QWDDf+zQr3hIbWPxj9t6nUXUsW1QbnFXYWgcLVPRv7R6T
z9wHuf9fHs1uR5oT0qb1wpkurBhifkiqLTOlcELf95dTBOhBajRr+LQYap1oiBvd
q/8So28EcRkgJbMotCYdVQiQ0NN9A6Kq9YWvwWr2vSg/5MHMGR4wfoy0743C1lXs
i2TE8BzZaTsXflr7CvmfyGttFikS2U12uuNT+aljsNt6PuFLZe5BZGGd3ocQ5KgI
qGRmRs7GXBVbsFhnpwLIrQI6h5rPthdoh2X3NW8Tok7E7QVj4QpJwiCQ/S0gkrEr
RjZYcBkOm0gu3wrhEwPv+mFPzEATQe3Ib1oLxG7hUi6VYygXsJDe51uhv9NF36et
RCYSWWl+lswX6s9iY8KNZWuTPAW+oefc30iAlaMdO/1bjdFfmbnZcnJ2deXPF6po
d/8ZodVh3EClGYTEaxJurevDYTz8HXQ5ll0CA9GnmT/SlihELyPAfjaeprW302Kp
aBQecU8WSCcMAYEjavlSsohhI11E6NR3xEx979EUG/gMSSLd+5aWFnTeu+ibdOym
42CCz1ju2amhJuHYKBnf8o4Un1bOkUcRV9eGnkAhlSe4i5vcCOR0xoGl20JZZYPx
GaI5en5p2oX6/9OvARgNJqgz2SYGvxT+6/3/O0ilOc5Sfq5JuihpoTqwjhqNsAYe
LZG4VAVBUh5yw/u4Vc9zdk/c/tEhJAwcD8mH680kcCHn5Y8GvQ4ThKDymv5w7ySH
gfkyp5sEpn0MuQ52mtyrfS6qmH9F6/ROUkZsjcYKFMmPDilAI0+xNcuuRJMEf0dY
UvfAHYHE4pr09eOO2S14meuKFS+6ZxxKKpqIC0A4NczGLTHaAdkSk4b4mLxAK5VJ
atfQFSXd5ymBjRIkpPQTKRHJSb0+NuKCXd3BIm0yIBKfND7x16fQYkWUTgsBnHhe
Gw/pvMOgEQRBPMajAWXnuVlUNNvawwBVpD+miIaLFIrSkKmTfaneCJDGx/veTNU9
S64ijmPp/Ht+mfufGw+F+BFOCeT7SVrlFQY9ea2AL0OLhZ296BKELfKd0b/PSe6q
ollZZA7Xu0eEa4xg8AYoy73byx5aUnU4sYU0y5jSQX7VfFF3Rbur+WlyMm47gnCP
CPfKPAbWom76ID5lsGynWkN7WoftHJz1j9PTz0q4k+jzjlUULvmP8e4LZkls7xK0
tmMQVo3rmWk1E4dq7Ek8mLqN3zl3s18HXIWGuXHypm2fZVF3H6QGIYWlcb4ZtMBQ
Wcg+HuzCU+gN2zRtJ4n7x5U7APrKiEo4zu4dJ6CHjX83wwJZjREvUt2yhpODe/44
myeFK/VoU3O63KdRMl2pqgmirs5dtc8obWxgjWIdAzWk8NchuZtNhVmXul5HZHb5
FhJihesLPCGsB3N9aiQ85hMgPrwdGHCFGCc1IyzHa9B1Q5K0YBD9Axd6L78/hbVR
SAVAANiippZdICu/vHeG2v0lRumRn7wuX3ofQVVJl+TVp8CajFgohAFnfBRjM65e
6cOm3Uqbl24H004WW3xAFGRuS/aAr0601T1o+EjMOEaRcXl+mr7XCl9i3bHb2l3Q
NHs5BdY2FcB1KTPHyZ1Ekh0uyeqt4CiVeO7uh5pWo2u6+VbL0lYZucf6kAEJWlcp
JR/6Fk/YQucGXSdJrvl1qScHWh5Gbbqm2PT6D9nktcsMO3z7go2l07Gl+kc4pGaU
zP+Be8bc9HrNxgvbk1tHv6LgJwpc2+7lH5M/2TwfYAflpUUUAFmuE9Y324FTMj0k
haPYy3aRhRHYNR3HOnh0nTbGSwFhrpxdrcA2JWyDZ5LgWPMYHbAXap+2QhdyHQ+P
GhmSCpiyi7AP0Hh7IAAuO5eAqWDanfFUaSTDJCT7v1470/bcFarNt4kTSpx7vRGO
UYMDbFx51xULNeiJAAbtEg8JfetYdB869jYsV78FDqgLStq3YEq3wxf9M4LNdMMd
XynaMw7h/TQGHQeKlhEYcMVwNwxvLihgLf5OezFOxIOizK4ViYEtFEKjyi18qhV5
mFN+5z6S85nO5Rxqsw69l9hNedsrBtBqr1MSSEo33CD5XPcj2K8CbnyabuvtXwII
1vg5M9j3Ixpaf1KG6AQC8WQRihXOXC/Jz9oSXjQCWQD/CVP/Qm7Sem8GiTO3b4n1
I+0Ka4nVdzd++MJ+e/9TfuFAQEAWPrUreNdOYzNLINhnrGKzwA3DlSR0A6VtphXG
zKjZXm7h10T9TKViVNMcfJXiSpTxl7aocbQmV6235dCvQT0Wa9MxUu3sJLlQvDYO
miff96n8vnJhYpM6bta8KPQnfKEIlNBo7sXhcI5pXnEkrjVWowJiSzZ5Mtg0lEgZ
t7QbBIiphQTJimfnNGDd3kkuEMhXpxu3b0JJx26sE/KLbsMuEmDTi5XKy6Qi4x9b
KRoz6KYKU4yfOdVRNLqCphY5ajarbC8yHCoXHyObFTZlxy94W7f5VroqxJjx0W6g
FsVTMR5n4IBLED7c8xUFSTa3RwyHWTSQdytVGonwY0R/mHlUv6qFA9Qqix9Ihc/f
J/WAaKa1yFUsveGBmw+2FXXaHWfpTILu90sxmHhAGl/64zdusQHH4hF5IJ1pH9ht
Aj65GJmx2VjKmAz66ZG5LATdYBYhPeLvdxXfLF8ZSJSTSHHhObF281Tj45bEcojv
SKrEFEOxcOwf0xSVK8mEVSi6hud47F2cIwdHTNWQlh1AjRSW0B51Qc5kk8TwJC2r
dfyDWXHY/HVUdUU1GD6V4uqrvLtK8aXr29QjSYwydbVeR46f0napi6JS4WgxKVZ/
42viluJDP67sZABiRtMLdgvnSrUc5q6CtKT75yR/xbTq/n43/NWVGlpfwy+rR14X
4zEv6PXrhkXDo/ofi5kgNFfb2JFK+j0jBi1OVOL9Qogho331Liaq/dzLYyH+QDy4
4BhWwP7PKvswKgksRsgkWyPxv9DOiv/hCL8SV42XfXgxI5qxt5ci9ACGD/WTF1Iu
s29/4ZJX88UiPucn295Nm9FiDB7fMfcA3KNft8v7hCNTRECrKqa84Z0yb4ZboXp2
fzBwelUMnzZb46hNxH944vZo+XHzVrC+Q7z/aMR4NAeIpPBilFLhMN4/XdJIYPsb
bQzKvPrYSARTqNLR1g6uT/yfp37itM39t1lVIqibmRqv2JN9co5dkqB1GCfAzYSO
ovlMc0Idwzfu6b+ueFcfNjPwG5D3Bmr64Ya4wIrezfxjXmzV5E6kRvrp43Q0x4m9
8SyaGa87Glu61gfDa7BsbygXiKMoV92SAGpz/66Ey7QHQx7YtHdiqbNzehfxaNzu
apo5NPsCVUbMw7X5EXG2wmvDIx6A4CpR6bhOOJNjawrx1O8o+J1T4EoFza5BZ2SN
DteEAM+1ysgeIyJ+kHA1oQlFiHtUH4KfDXaFha3nEO2ea8ktGXGsJayOZeA2520i
5PvipKTwt0nkWTuOgU4Wi6rxlLeS5vr+lD1Ttj4yrJQ=
`pragma protect end_protected
