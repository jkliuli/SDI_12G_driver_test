// sdi_tx_sys.v

// Generated using ACDS version 22.2 94

`timescale 1 ps / 1 ps
module sdi_tx_sys (
		input  wire         tx_core_rst_in_reset_reset,                  //          tx_core_rst_in_reset.reset
		output wire [0:0]   tx_phy_tx_cal_busy_tx_cal_busy,              //            tx_phy_tx_cal_busy.tx_cal_busy
		input  wire [0:0]   tx_phy_tx_serial_clk0_clk,                   //         tx_phy_tx_serial_clk0.clk
		output wire [0:0]   tx_phy_tx_serial_data_tx_serial_data,        //         tx_phy_tx_serial_data.tx_serial_data
		output wire [0:0]   tx_phy_tx_clkout_clk,                        //              tx_phy_tx_clkout.clk
		input  wire [127:0] tx_phy_tx_parallel_data_tx_parallel_data,    //       tx_phy_tx_parallel_data.tx_parallel_data
		input  wire [17:0]  tx_phy_tx_control_tx_control,                //             tx_phy_tx_control.tx_control
		input  wire [0:0]   tx_phy_tx_enh_data_valid_tx_enh_data_valid,  //      tx_phy_tx_enh_data_valid.tx_enh_data_valid
		input  wire         tx_phy_reset_in_reset_reset,                 //         tx_phy_reset_in_reset.reset
		output wire [0:0]   tx_phy_rst_ctrl_pll_powerdown_pll_powerdown, // tx_phy_rst_ctrl_pll_powerdown.pll_powerdown
		output wire [0:0]   tx_phy_rst_ctrl_tx_ready_tx_ready,           //      tx_phy_rst_ctrl_tx_ready.tx_ready
		input  wire [0:0]   tx_phy_rst_ctrl_pll_locked_pll_locked,       //    tx_phy_rst_ctrl_pll_locked.pll_locked
		input  wire [0:0]   tx_phy_rst_ctrl_pll_select_pll_select,       //    tx_phy_rst_ctrl_pll_select.pll_select
		input  wire [0:0]   tx_phy_rst_ctrl_tx_cal_busy_tx_cal_busy,     //   tx_phy_rst_ctrl_tx_cal_busy.tx_cal_busy
		input  wire         tx_phy_rst_ctrl_clk_in_clk_clk,              //    tx_phy_rst_ctrl_clk_in_clk.clk
		input  wire         tx_sdi_tx_datain_valid_export,               //        tx_sdi_tx_datain_valid.export
		input  wire         tx_sdi_tx_trs_export,                        //                 tx_sdi_tx_trs.export
		input  wire [2:0]   tx_sdi_tx_std_export,                        //                 tx_sdi_tx_std.export
		input  wire         tx_sdi_tx_enable_ln_export,                  //           tx_sdi_tx_enable_ln.export
		input  wire         tx_sdi_tx_enable_crc_export,                 //          tx_sdi_tx_enable_crc.export
		input  wire [79:0]  tx_sdi_tx_datain_export,                     //              tx_sdi_tx_datain.export
		input  wire [43:0]  tx_sdi_tx_ln_export,                         //                  tx_sdi_tx_ln.export
		input  wire [43:0]  tx_sdi_tx_ln_b_export,                       //                tx_sdi_tx_ln_b.export
		output wire         tx_sdi_tx_dataout_valid_export,              //       tx_sdi_tx_dataout_valid.export
		output wire [79:0]  tx_sdi_tx_dataout_tx_parallel_data,          //             tx_sdi_tx_dataout.tx_parallel_data
		output wire         tx_sdi_clkout_out_clk_clk                    //         tx_sdi_clkout_out_clk.clk
	);

	wire        tx_phy_rst_ctrl_clk_out_clk_clk;                 // tx_phy_rst_ctrl_clk:out_clk -> [rst_controller:clk, tx_phy_reset_0:clk, tx_phy_rst_ctrl:clock]
	wire  [0:0] tx_phy_tx_pma_div_clkout_clk;                    // tx_phy:tx_pma_div_clkout -> [tx_phy:tx_coreclkin, tx_sdi:tx_pclk, tx_sdi_clkout:in_clk]
	wire  [0:0] tx_phy_rst_ctrl_tx_analogreset_tx_analogreset;   // tx_phy_rst_ctrl:tx_analogreset -> tx_phy:tx_analogreset
	wire  [0:0] tx_phy_rst_ctrl_tx_digitalreset_tx_digitalreset; // tx_phy_rst_ctrl:tx_digitalreset -> tx_phy:tx_digitalreset
	wire        tx_phy_reset_0_out_reset_reset;                  // tx_phy_reset_0:out_reset -> tx_phy_rst_ctrl:reset
	wire        tx_core_rst_out_reset_reset;                     // tx_core_rst:out_reset -> tx_sdi:tx_rst
	wire        rst_controller_reset_out_reset;                  // rst_controller:reset_out -> tx_phy_reset_0:in_reset
	wire        tx_phy_reset_out_reset_reset;                    // tx_phy_reset:out_reset -> rst_controller:reset_in0

	sdi_tx_sys_tx_core_rst tx_core_rst (
		.in_reset  (tx_core_rst_in_reset_reset),  //   input,  width = 1,  in_reset.reset
		.out_reset (tx_core_rst_out_reset_reset)  //  output,  width = 1, out_reset.reset
	);

	sdi_tx_sys_tx_phy tx_phy (
		.tx_analogreset    (tx_phy_rst_ctrl_tx_analogreset_tx_analogreset),   //   input,    width = 1,    tx_analogreset.tx_analogreset
		.tx_digitalreset   (tx_phy_rst_ctrl_tx_digitalreset_tx_digitalreset), //   input,    width = 1,   tx_digitalreset.tx_digitalreset
		.tx_cal_busy       (tx_phy_tx_cal_busy_tx_cal_busy),                  //  output,    width = 1,       tx_cal_busy.tx_cal_busy
		.tx_serial_clk0    (tx_phy_tx_serial_clk0_clk),                       //   input,    width = 1,    tx_serial_clk0.clk
		.tx_serial_data    (tx_phy_tx_serial_data_tx_serial_data),            //  output,    width = 1,    tx_serial_data.tx_serial_data
		.tx_coreclkin      (tx_phy_tx_pma_div_clkout_clk),                    //   input,    width = 1,      tx_coreclkin.clk
		.tx_clkout         (tx_phy_tx_clkout_clk),                            //  output,    width = 1,         tx_clkout.clk
		.tx_pma_div_clkout (tx_phy_tx_pma_div_clkout_clk),                    //  output,    width = 1, tx_pma_div_clkout.clk
		.tx_parallel_data  (tx_phy_tx_parallel_data_tx_parallel_data),        //   input,  width = 128,  tx_parallel_data.tx_parallel_data
		.tx_control        (tx_phy_tx_control_tx_control),                    //   input,   width = 18,        tx_control.tx_control
		.tx_enh_data_valid (tx_phy_tx_enh_data_valid_tx_enh_data_valid)       //   input,    width = 1, tx_enh_data_valid.tx_enh_data_valid
	);

	sdi_tx_sys_tx_phy_reset tx_phy_reset (
		.in_reset  (tx_phy_reset_in_reset_reset),  //   input,  width = 1,  in_reset.reset
		.out_reset (tx_phy_reset_out_reset_reset)  //  output,  width = 1, out_reset.reset
	);

	sdi_tx_sys_tx_phy_reset_0 tx_phy_reset_0 (
		.clk       (tx_phy_rst_ctrl_clk_out_clk_clk), //   input,  width = 1,       clk.clk
		.in_reset  (rst_controller_reset_out_reset),  //   input,  width = 1,  in_reset.reset
		.out_reset (tx_phy_reset_0_out_reset_reset)   //  output,  width = 1, out_reset.reset
	);

	sdi_tx_sys_tx_phy_rst_ctrl tx_phy_rst_ctrl (
		.clock           (tx_phy_rst_ctrl_clk_out_clk_clk),                 //   input,  width = 1,           clock.clk
		.reset           (tx_phy_reset_0_out_reset_reset),                  //   input,  width = 1,           reset.reset
		.pll_powerdown   (tx_phy_rst_ctrl_pll_powerdown_pll_powerdown),     //  output,  width = 1,   pll_powerdown.pll_powerdown
		.tx_analogreset  (tx_phy_rst_ctrl_tx_analogreset_tx_analogreset),   //  output,  width = 1,  tx_analogreset.tx_analogreset
		.tx_digitalreset (tx_phy_rst_ctrl_tx_digitalreset_tx_digitalreset), //  output,  width = 1, tx_digitalreset.tx_digitalreset
		.tx_ready        (tx_phy_rst_ctrl_tx_ready_tx_ready),               //  output,  width = 1,        tx_ready.tx_ready
		.pll_locked      (tx_phy_rst_ctrl_pll_locked_pll_locked),           //   input,  width = 1,      pll_locked.pll_locked
		.pll_select      (tx_phy_rst_ctrl_pll_select_pll_select),           //   input,  width = 1,      pll_select.pll_select
		.tx_cal_busy     (tx_phy_rst_ctrl_tx_cal_busy_tx_cal_busy)          //   input,  width = 1,     tx_cal_busy.tx_cal_busy
	);

	sdi_tx_sys_tx_phy_rst_ctrl_clk tx_phy_rst_ctrl_clk (
		.in_clk  (tx_phy_rst_ctrl_clk_in_clk_clk),  //   input,  width = 1,  in_clk.clk
		.out_clk (tx_phy_rst_ctrl_clk_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	sdi_tx_sys_tx_sdi tx_sdi (
		.tx_rst           (tx_core_rst_out_reset_reset),        //   input,   width = 1,           tx_rst.reset
		.tx_datain_valid  (tx_sdi_tx_datain_valid_export),      //   input,   width = 1,  tx_datain_valid.export
		.tx_trs           (tx_sdi_tx_trs_export),               //   input,   width = 1,           tx_trs.export
		.tx_std           (tx_sdi_tx_std_export),               //   input,   width = 3,           tx_std.export
		.tx_enable_ln     (tx_sdi_tx_enable_ln_export),         //   input,   width = 1,     tx_enable_ln.export
		.tx_enable_crc    (tx_sdi_tx_enable_crc_export),        //   input,   width = 1,    tx_enable_crc.export
		.tx_datain        (tx_sdi_tx_datain_export),            //   input,  width = 80,        tx_datain.export
		.tx_ln            (tx_sdi_tx_ln_export),                //   input,  width = 44,            tx_ln.export
		.tx_ln_b          (tx_sdi_tx_ln_b_export),              //   input,  width = 44,          tx_ln_b.export
		.tx_dataout_valid (tx_sdi_tx_dataout_valid_export),     //  output,   width = 1, tx_dataout_valid.export
		.tx_dataout       (tx_sdi_tx_dataout_tx_parallel_data), //  output,  width = 80,       tx_dataout.tx_parallel_data
		.tx_pclk          (tx_phy_tx_pma_div_clkout_clk)        //   input,   width = 1,          tx_pclk.clk
	);

	sdi_tx_sys_tx_sdi_clkout tx_sdi_clkout (
		.in_clk  (tx_phy_tx_pma_div_clkout_clk), //   input,  width = 1,  in_clk.clk
		.out_clk (tx_sdi_clkout_out_clk_clk)     //  output,  width = 1, out_clk.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (tx_phy_reset_out_reset_reset),    //   input,  width = 1, reset_in0.reset
		.clk            (tx_phy_rst_ctrl_clk_out_clk_clk), //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset),  //  output,  width = 1, reset_out.reset
		.reset_req      (),                                // (terminated),                       
		.reset_req_in0  (1'b0),                            // (terminated),                       
		.reset_in1      (1'b0),                            // (terminated),                       
		.reset_req_in1  (1'b0),                            // (terminated),                       
		.reset_in2      (1'b0),                            // (terminated),                       
		.reset_req_in2  (1'b0),                            // (terminated),                       
		.reset_in3      (1'b0),                            // (terminated),                       
		.reset_req_in3  (1'b0),                            // (terminated),                       
		.reset_in4      (1'b0),                            // (terminated),                       
		.reset_req_in4  (1'b0),                            // (terminated),                       
		.reset_in5      (1'b0),                            // (terminated),                       
		.reset_req_in5  (1'b0),                            // (terminated),                       
		.reset_in6      (1'b0),                            // (terminated),                       
		.reset_req_in6  (1'b0),                            // (terminated),                       
		.reset_in7      (1'b0),                            // (terminated),                       
		.reset_req_in7  (1'b0),                            // (terminated),                       
		.reset_in8      (1'b0),                            // (terminated),                       
		.reset_req_in8  (1'b0),                            // (terminated),                       
		.reset_in9      (1'b0),                            // (terminated),                       
		.reset_req_in9  (1'b0),                            // (terminated),                       
		.reset_in10     (1'b0),                            // (terminated),                       
		.reset_req_in10 (1'b0),                            // (terminated),                       
		.reset_in11     (1'b0),                            // (terminated),                       
		.reset_req_in11 (1'b0),                            // (terminated),                       
		.reset_in12     (1'b0),                            // (terminated),                       
		.reset_req_in12 (1'b0),                            // (terminated),                       
		.reset_in13     (1'b0),                            // (terminated),                       
		.reset_req_in13 (1'b0),                            // (terminated),                       
		.reset_in14     (1'b0),                            // (terminated),                       
		.reset_req_in14 (1'b0),                            // (terminated),                       
		.reset_in15     (1'b0),                            // (terminated),                       
		.reset_req_in15 (1'b0)                             // (terminated),                       
	);

endmodule
