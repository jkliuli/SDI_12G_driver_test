module clkctrl (
		input  wire  inclk,  //  inclk.clk
		output wire  outclk  // outclk.clk
	);
endmodule

