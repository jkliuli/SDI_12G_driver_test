module clk_io (
		input  wire  inclk,  //  inclk.clk
		output wire  outclk  // outclk.clk
	);
endmodule

